-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dsSq/7wK2XqTt2Uw9VCuhO4oSt5kUlQFu65wLTBbdPS7dhGRXJH78rnXHTpmeMlyz/A+RqbjfCKu
HpZ35TpHGwlwCKKTaXDGGxqBN7bWJ7toyQ17S/m+9jwMz28iOiP8hgZw/X4FD5RJnSAkeu9vVSKB
vhEAIha/fNwGesbMUUqA3QcHnV55xcWwYY39zSd4jFw+Rl7dXDq9J9LPcunWE5z28QQjI8J40GsM
Zl94jEVxEafPnyK4JM38MFSKyideZ/H5RvmYezdjZ6epizZhZIVVvveGmO0f/jipl9gkh8Kavw1P
0dGQQkz+tWRUq9o/qIOgyGE6u25c4cAERx3l7Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25264)
`protect data_block
uXXqkRuF2n6jnIcSNfxBD1vCMyU03a02mC3UBnJUehT/zfUmY2+r18GNBE5v5M28fZE9x9WmZRcd
Dk54SdKPfU6UGyGyCTtN/Oa09RdaL33BIPJXVsXFIK6g/M+k1aJB9yteM4wVSiZM3klVMImQG4hL
+Eyu4QrzmmcrvCc2uDWGsschzrNPGe1uMesT/gZ2ovQ0yWCKQgjDNFPSPtQT6aBnUGyYKW4lD39f
KUJGTCY8gIwlQcBAd/Q1r0OKYuwKLM9B+Xd/4rq632YHDntyoQrLlIgZZSjfueyJJVaVXh0kD6lk
g9AwXWcH3yb1q8ehBpqBrjNV/NiPdgtOb+7mRaKRD8NxnxQ8y0YDRx6ODTHIQktLCB/Od24j/CtI
MzB0XYZKVX36KboCHXpV8kJ5gi88qplR7nDx+04hZSQurNCavWu93h7433VJmHYpC7Vtrw9kDmFY
ZpdQx+2uM809m2V4lg/668XTHp1aVejqpVTOkpiX3VNJgHUqr8D8O0fMNsoT+d/1zslflA5k1Dqs
0b3c0IctMSsfLxQOP52LlcziTbLoHtjuT5k+lTVpGQ07cVKmZnbNkCXM2yiV8ZQoIWYMNsAQ/oH3
HJFS3fNgqVBJnSMHO273/DL5s3zLLjKeOvBK3vK8RA8NzbVNvhvuAIANSrtjdIl8fJ34A1V3QZ0t
UHr+SbOHUWqAPrZQckeoePJx5va70y/OnoLp+pmQouSo+ROf8OJSwg399SE/LS911cCml4gDvSM2
DNblRGBlFTK+UaXS4l2jgP/72kCQPWzs7N5juwz5JQ/0gl0UXNlG7p6meS8Xg0y73k8a6PFmSysk
HszXBhaizS6pcmuQFg6DUzp3DxtPxuU0BZAgj564udpldE5X3R6oxRKMAaddyO2ar34n4EJwF7s9
Fud796voDTNboqaD99PuDZtxB0s+ux7xffjNGS0v+6dBoepGGzFV+pbos/cqQD9W5vrDa0T9A1Lk
kt6VwGhsYyeUBraWBPoktmLRONX32t2+HUh4B9lr5abw77fOEaZUz9EghjekB0xeD8nYv+SBkZfW
Bf6BIbgRPobR63xCsPJmjJe0USDnxaSNS55h/3tAfMAyCwU0uF1G36iIRwwH2s8gT8Zag9DkOkU0
xrqP0ofpxC4csAFaU5oirKfGvkmVNyFNPjIbuYVo7nydhFG+J9xbdd7DTZtJ9CdrBRztxaVV29Ec
/ndVqMEuGBPCqpzbdqsX2vBvxgHYG9djS08UhG1t+xJWn3LUdjssbpKxp9iykgNSs5FmZaKnpLny
eUAMD2Hhx0h28+nr8TF1PcDJ3cjxUQFq/VBLTnz/4EaFYjN5Cho1hOKcaXa2mqkVLupxDWnYQ5vJ
kTWV6tBcaExCqOFWDGwnRAz7ULXApKNr6otg+MXZoDma+83hWJAWRFpIwccrnqdD38zLWdd1n5W3
3mmMqO1dQmYcfrIpt9gdQWRNWvYLXSB4T9el9mriXbSjEkC/XbA1IR+Zo5ugZbHMTus0PNZYvbM3
C9dULvQL9xoxmjdII14Fn9DZ7wLRx1s+Vt7l0CwZZ4iZ22S7dNFGn0IIvMW6oJ/N4kUKpDDo+clf
DW2+cOwzN9KVZV7VYaRGgYzkb76nnFbdJ7shK5EcJdFIdPEgDg0LT6YtTx9G2zUFjJp69L5DYKos
xAhg2Ml2orENXICwdnaKTeJP4H3M8ffZx5BwFKb0oULLjdb7X4CPRqmmMfv6zhk9MODX07rqmUvi
SexQOgFL6Eh2HGsbafsdbw0+5mbldlPuuUmZFRGe5J1nAEUQo0LpPD398/rnRd+q2BcP3eTNf2Dk
8NJnw2jRN5u7uDF5S9fgTkwdKqHr+CjqsiNw85sgXltedxzZF3qUDq+N8fr/xp2/1o/0aOZgKtgx
YzLcjdw9OaKU1UFliSF9KLdNEGmpuaxTeLsA+wa5rfT9wjd4c3UeBlLMypreg684w+86cNN4EIHv
ONv7fiLrGfo/BRgbI9JIGnIdITph5hdDUDCrk2YRv78Wu6zvLYp7YEuuYV6peEPbnWWA0dkR8JwN
OvLj6LReKpoxL68sNrHJ5Go2etdf/jiOz0NdIC32URn1bCWn2wFbcmY+iNeK7SVg1ZJyic39qj7N
/X0aFye1Jt7u/aNOBt+AWX/YJ91AU3k/cwVxb0O/lbfCjsvj2zju6mBGNg5t6gJEAax+14WERqZm
gcEqPiiJOUS/OYNYnZpPmCnt+ejGYJ7kPWqEW8WOP0KSxuH+BlT5ZRD5hNnyXU6BUmGIBpFHCb3M
+bYJhx4Y1VXEevTuQzlgPaFZMjWlnGfmAl7oXOtMiILSVxCqP6ElW55rSOxqI+VHGJsetzJOhRBW
iUGOB0kYbkE9Db82psd6cJRUvstwyeL5rAsN7gY/rYvIUVnIr5o8p9bJa9vxYqotdNd3AYSd7AD6
eocJoHelPMAh0VJ9wh+xfvw89mezGJounsbDU66GKlqFVtSLewlafu6GC481rVabFwWACLHYa9no
CNNWpcPEtgVhDM6Dc42+ZICClkGYQNnfQzM6+ihsmsa/hcE1gKLwtD2XdHSJ8tuoS+S2MltmMAlz
zKZAA/jyD/UQ1kx/8Y/KgBPDQB3zJrrbTXf9IxOygGqYsbuYDFkM8RDucAFG3jzzB2y7So7yVVv8
Eu58LasHwmThdh20NFr2vEseASKmXIj9Ib1HlkoUMZrEeFj0AOXaQ+niJffTqyTE1dVI5a3ZKrHd
a/WTuLtWgsILCdFjK281X4vWMtcA4GEacESRfPEvhdbyaqjtlkC8zJhMVARBzFar9fitppkXWDXX
40i0wCDICBujsYbM6/88FjnvYWEOH8icB76qWrQ2UBruRm6RnPIFkuJS/E90McCJCvh/nInGZ4TK
j6p6+UcDDzg02vm7cz+cSbEtEphqh9jLBpoU8v4hHRkxzWHJFcNojCeCJGMlEdvazkUCFcO3c9xJ
gY4TWzK60pSpgoiB8GEuNNiePf1G9EWyDtA9F8PfqRn3wBfiRuPLCJJ4440iKMqgfUQlDEThMPGi
BfSQ6e9S+XvJXwBHZ0ATHkosL+rf7lBV89l5ocbdyH2OWig+Pt7pM576qaO6Z+xaJVTq9SUlHC8D
tavt9jtHp2GuqpQHeicol9tb/M+6ojf4QsLcxmQ8wUh+2fvcvev5aTd6m9/OyFbE9g3gmx5tnWiR
CBUn+ZXpJPGGCkQePTSRw4jLCSQ5Pe0+wj0dFunLKxpPPKmtgm5wUMUGsa9LrzmO5czV5D+jJHZy
s7Te+rjxq7wA0Fw2t5ydNiCZR03m/yyazprCvTmHwGsgK2/eI5wI2QBPQ7uDG3WSzJRk5qYbTKON
2sVOGeSdnYX+oJUCHWDR+/8oBLT02Gmgkh0T9atJgtT1ZiYGxEmqau4KT1tRieJTK3GA0z/li+Vd
5SOBYCgJZKpghPTcpNWVXz/71EGeT1WUlKJJpHIMudjchv8bGq/BTGjx6RmCYCcjrCs9q7WEkdjZ
gvVJI/Ow4kcE0OBm8RQz4RPDkU03AmfucbAvfFpy7WWN2QTFGr1x6ZNW7qe4qiESWBzvPB6TveJq
CowBr2rvSx56jU8evfQF01vww8LiUipx5opnstnO1f86JCnymK2e02nBAXaaZsOoBU0eQRfFML0L
WZ1Eu0828EW+5H3w1lMqe7EwaJSHqCHVgoWPmXrID+BMgeX6luGKEtSlLevr6KUk/iHItaj7pPop
x1zedYMlUr4bQk1rdglRamOrskkpejKASI56tj4toAS6/z6WzrulCe2j/ltaXip+Po6HMmX3rPoC
seWa/ih/o800Gx/wex83PgjHJdgku9FmYLdjI2v60cf3B6wU9QLjpmUUnaCL85Sr8uR5hYXhC3Tr
B/Qu5v2yyCUe1YNy15Z9IMHqfsCJdamNCJ7msB5xYB364fcSsubAsQ5wVNH4PsVRenLE/3gRydCJ
ckRPmPDd0VjBh5Ai3AhSgaMuY49itDR/u2sMYeBhkxajVfNoytbunhmgQXElXzQfORCcDP7xzrdp
RJAnWvDAhvIGrw6NERHsctrwWnj+ZWxtsl7rfLyZxl2kmsvtWGN4WjACq0tzCXsFeDrI2Ysgn313
6llL2tEvTjgU/e/7f3pQtboyA9bHUJhnISwaydmLYZkmZqfNv/sWBimM8McBWipgGLe1XB3n8rmp
DNVX06UYtfHsmyrLWVOMxNnc982h+moLWdre25gBLS8AmlqxkZmXqnF4+usQ8WHfDJSJsf1+gUML
zcHWGaE8pCQx0kaz+KpsdFKUyKXzHcvSLORfExvtlyIQN3KjqWFMZY32EtjO9S4hhNkldxTS9j+p
mh3Fir1aU8HL3S4bvC9IcJ8ftxaU2UwmCwcOT1jDJMVR7ku53eCkj+ZwgTK+jx/kK8rYdTsq0gky
ka1FFM5L0xfMcvKOJjrA/yknyEnAqZ70AB8ILWIZiqnUEdBnsZYxKT/ZGbfaLBfxbavc9PkAwr1C
60R1RvGeBdw1NQWHphyQl1iMoM0oW1j3/PWzsjhhTj3hJK3pu4KcvcU2hVFvywmmrmEJEAxm6dyi
ncg8Ow4Mpvxe7jXLvuxLZEBrSGh4+KNgJLhYkqNBQnlN5hmQLhtxCdzaX91dN92IiyByc5ME+c72
tResgSAcZmcLKDDldaNrBMOYJ1uxLwp5DdqCxslvpK0leFahtYbHWQp+I88+VSEhAFScVsXB5tIS
5Inu1VDT8iE+H5aW4mgMj2waE3tGnahpuvzacgo2GPVEmx17Dh3rlExCZNyA6cwS9zA0JuTUPhP7
Kt7eqS8HkMJ9pnuAwDDA7kmfF1eLjoOaDVUk/M6lxUFlFH49usjX/vTnf3VAS2FnarwEcHK1Y93r
mQfADhbwCdO7kEpGIaYc1X37fthWNuODC/bMxKmidJxVUi1il6cKgto49YMEinEKDDxiZWEKPjWH
6g2jYJnuyzXO6nOGwUad/e34Seaf5NgvjfRW4Xz7WhShBw4iPuBRg0Bogzg2J4EBe2TVODlxYT6I
VE8SD/mDUgNaG+1bH5gLI1OZBrA8X1Vbkc9d2d7PPWoLYMyG8p2vMKeuS7sVoA/xit0wt1r0X6Do
aUJc7mMk9N83+VJT/4O2YbfzSSuY0ULuNAYhBYNU1FLbrhqAd7YpsSJa9xstolrdovklRMKxg0Bb
7qMSMKQ8lTek6CPXou/kTnzVkwssKlprGODUXIeeDl4jB+NR3ze+uhiwG8js8DwNB9t+Pg//+y3r
wR8fwvHpy+/wAn4ZepW5Mg4XL1ZjYq0Mp1iAEAXY6UXdXocrbFfhMh1FDQwL3jNEiW0d4ONahmpV
rCQUDMPUscmDi8noi51jdt2urSJ/lHFQU+Rp+uqac8pOtenqa9n6Yql7APOaRYDi3antIEFtuUnd
TzE4frguInMic2HG46Oh11If8Tyn5FcNrA59lpq9+otSHoTePhQjyAYctCDPWymtIiRp1ScIwCTV
bVzvBZYB4blQ1YNH9PQjsSYOWxPRAKpEKzXAP1y2v2mirs6JX7s2mJpi4m5OX3uklIYYaSrNHjKF
sM62mvb2sdHjJ5VY4H/73l0aoMtGWSpUjlo5ATfxHdEmvnDJciawfUgjeBy4xfmkaT4UCDy6QqAk
k9xJerVgBLs2uEDNiqAg1CPVR7qr3Vy7DY4OMgns6fwwLDvG6ebtmqbJNhpw28U70jWri6UKjNzF
wLBnZXsRHaNSwa1BBhp51X0B7Tkrvry6iaKVTS+cjrICQqWemfqgJRfamXEftdLA+IkDhF49XxcZ
JqwyrFMvHY1YZsEK92XBG1svbNx6zs4x4KaNslkGfBhZ8ZFhPWnELOoipJRSIrhPllP3cgk/cm6W
o4OO1MBahhl/ZCyTs04w7LiiOsgSMFbx4lC2odMvblOm3uEMACyt+6QACAh35bmtk3eLE3pOJm3L
Y6c8JtR9nJVOSdRtAV/rN7hOZfTQnm7QM2w465uUKbnOxLuXuYLFWRWnHyJpY5pCwFaYaJntzw8H
M52urbGrretrDYgxr1oyLnl8kZ64WAVrm1i+NTJkFNUqOv8qLUj1ukGqU/gH3Hs97+tqYRsieg+0
kfmesZMNh3h6QmORKcJFi30SDn/llqZBZq+uyrqyf4mBLpdT4NBjV6bw2rAWL36YmROG9WVb1L/X
bZMoMh7cWp+AadTyxDR/YaAhPNa9w/+PSvOzId3C0V9VrzBQ88OKPPK4diJyYpFTRqP0Zi4vZIzI
Mq4zJN9IsMbGx0UMlVn7gOvp2t+13ohgQ9ThlKoS5mSNKsB2j2YxPRcWcEn84ydTClP9S91W022g
JwYZYHnJwsO/Z4uSb5jBMhgIeOSvuvFRuQQF69VSrVpbGRRdwMYnCGC5fH8urT4RmMSie7/jVj2F
FwR6yf/Sf5p54EFo3NCoiiLXCfyMymCyh0Db/YSAlMKOvWgF9DWfTpUoLfgtTmn3CwSBXEYO8wxx
R8E+MIfP/9dAw8gy5Q/CmwSFuiWeFuUGkVZPgZ/xSLTeaXE0x3T3ChIeQGvqR84pecb4Zl9aYQLA
H6BHCmR+ybSRp3AgHxKPYGF22vo5FF4DXvoUwEMsSS6gemXkbasxwYtjDj2YfuCTfTOFvVRbVHut
cz4YDCdcJzMS8k0vxo2lMJChwP08+NVXjfqAPRH+pqXBkC2LJdIwzPWgCm+p3sSuScpfcCH1Mhjn
8AYq/jnYTcJ8TUrGpkrLeJ14z3aMZlNKJoVfBFcYXZ/1L91ERUrGB8+d7GC83yyVfKfj4i8GREV0
JryVUOUAuOeOGbNitNw2VKybmT6kW4wyTai+2BL9Bku0uzXyTIGUFQiOnjGp1B173fJi7UBGIC1o
TCN72ymHONp8AdjE4x/pSNsq7grDhEU6lVl0thOdTVrBU+GCJQ1I3VlCvaH8C18ISA2bdZLZGUdT
73gkgZMMef40Jmr61V7y78wUGOmCYoKyYwV8lMNUWDpamlgH+aWA+0p2ZV+7BGP/cCG5OoHVyG4Z
73Yjm7rct3v8J4FhTeBY2w9xcg/7QkoApgQt2wz5pStkgzCGkavCU0ljuG3Du0ASw+fvWTm7gj0F
KiZoNPJzx2GDozeO5P8hjT7NzEQ1tY2QFEnmmgBqmgQ4VycqIv/MBaxpzVt4W+GuRgzp0Yq5dRkw
QDNJLbPkOHemiCvn5FVSCTmqytk+IbQ/QKyUq90lTY+vT/+/I61PU0dFxtSORXl/J68XaA2tTxfW
h1nlQhLvSQl9j+V6JvZ9l4YW5tc8xI++yg0Qj5InLmr05GppR6Q+ElhtVPF/SWzlf/etBUgFwXS5
JYJy8YgbwVNZMtlrPmWEApQzf2NMCRFabDGud2ZowkxRVIjUn440uN+foHmXFscVe4NemuRODRFY
EmV5+HSdkqN7yY7vAxtgFDCxHAex8p+Fr3PlgX+QkjGmRdQ7V9aDUICIzN0Li5FhZF5GvKS6DVK4
WWZGDuG2GQ/hFxoFDyMmCUxP5QfCaf9S7NemUmagxKdXSLVMUUYOJ4VUYUDIKHGIaYiSuh+MgG3s
eGxCVXSC5qLXgSB9ApAkvYUHvGlu44DmZS7qbqdphCO6E5MuI0rpaU22jKQKgFPLPq/XfKzjfNQx
xLkxSjbEpihQRGbV6isdhgOckyrdeoQJEPlkiFfVHAOtzjoO54hx//auQbwIIdsH4kWphzmmZImD
xM1dskumtVR+9KjWB0BOGXR2RTPPlXpQiw/+kr5EddBe1U4Ezeu3zOLLUy5DOcQJ3j6vo7/6ktBw
WZP+7LjD9qP2R0O1pf4Uc+xc0vfnioqDnrYlbodRD1wWEgdtUOAoFoLoElrfZGVmx+WXRkYP5+dD
ucCk6zmkIU5MnLHunTevsYTlPKKstfJxDX0fhMbq69aVNKpcw3Cqntawyzv73WDLm2/dxntt9j4p
aGhh6NclGjuKQ69wxCZ98YDe0p5rON4ikKV5aFLZ/3JHZgDTHGRXRkyy8Iw7zDydNsdPmSiKpsL1
ZsFgXtCoKaGgjiuo+QcluECx2WTCl6GcUnnNAY40upjlX0hVUw4D9j3Pzz6HbhvXANe3up7w4JTv
YKNIrAtYZlJ4Cf+YPOajl+XEl8DvNjViAyaToz/v5JyYFmijfE5i07LlIgMiiSSRw7WPoqCtaO1a
gtd9ESrsreGWkErsOqyXE2q+emm1tDz0oRRX/bXxCWA1OrHutl+B6UlLU5jGHak5DyfbxUPngiQQ
RzZbLMxXl/RPTTvEKoPSpNKNCGpF6ayTHfmN/pgmW71G6LLB0uv5LKjrXyjopPu0SNCCtOqvWt1D
Ma/ta7uHiguuXoaD5RhU51WnhhTuV+z2ysV7YUVZ9lPlefNGfaJOBAP97A0T6vzUHXdNFOkxhLma
fXVxu9OFUug/Z2ranUkUq8Dbro1rpTZwAHXFYnsQIWe+NBK5n05J8+iVB65F8ZyhL0ntCvbau1z+
y+QHpO27FZltXg1qhEjt+rs3kxzcCOjVK0MEB16kkpRGwvsjEqYX02LCeVwjUQrC2hdMDobNMrHg
0KNjTr+t8pElOfuAKS4C9AEH5MMtMU/m38NC603HL24NlQNwPY4RVsRVCq3+hF1la2Zqn7Mpp9QR
KZJMsOffy8QfDtIccP2h+N2HFR+J8senCHvLoF3sOEj8yRqqSGeC7mGdeHupcCZ0C4wGz0BJvv7Z
lP3TzNZRwnJ+rrUfQQUrKTqoEDUHVU92OS1yrWa92JbJV2yR9Wo5KrqRgoQJnvZLJLQz+p/RzeSC
SKujkrpbFRALvyKzMRpF3Y5icE4eUNB88VrjZprjms0DsWiv5cRWLFPYmSpkaz1eVKTEsTmwA6A2
tm7WwBF8cIazhIY0MM+GtWI38ulw022yL5j7xeXuzJGMVuytBTAoaW3et+rtKcZiN6u4Aob3WkHZ
imm8ZfvcMOcw00ye2qDfyOfo4mcfVPxpI1xLmkdGwAA8n/fh09S36jxUp8W1+YOlN/fAMLmzb81Q
gTtQQoD4uptR7ocsu+fGQpamCMer13fWAuqt48kElS5O2J0inii15etyZbW3Hh174YM26kR0Ikkr
ZXjN9CclZbaGkhFx94mNo+XEq8TE9pq2IU88gm0OEYmFeQKbLf2LG8p5bTgaMUZlTOOb0FFjylRf
a47kJEaQtwRA8Tj0CWe8pE93e/0CsO2yGmy2txCSRJviTQjX+9PtUeAff6bc851ySvsAZOf0N0Kh
5TNy6VqT/n+lsNNBIMepKRnSGi+GHunrK/Jx+9KCierR6IiK2/VevpOzuS1cWAWUku6GCjyHXpN9
0059skYeCxCBy+gY64VLI6uergqPFcccGySCNqiYjdAMFLrQtTRJU6vgZVQatWHnZuW60VSid1Ef
apDOUnUPazL20fhO+xogUIyRJTZKScYJUzYUqU9X/zqvK+tWTR0t1fST28DKQO+LVaJhyrhyOtTL
HFDzxuRVDrv3Emk/QSgmX6O6w0fWBwb1cLFj7v14CpVKM2vvonr1ttys22MJDZR5W700HLur0FGU
hUdSHxO5zRlhdn/tJo6y3YvEP3/ugB/PFruoxc9T4kTrOmAtuv3RUfKXG77zVsncJikO5z/c8IbH
NLSexG5fMqaVC9k8RfER2qWk25lu/IqRvdmHnUKD+OQcTbRz+XeELSyG+ymSauz5fBE2TMtzXmAf
snVA9yqH2Dq54MJF9/DIZtCMcPq5YMQ0xep31+oBfq8K+8ZNeaNPoktze0UQf3bFobRaqosaggQt
UqIAhe+Mblmkc7tEeTQ0ZWFPdkBL6AlYqn1XRCvNQ0t/HqOsmJGiiWwym/Na04UxGSyRjNke36Ck
nWOaI0YquMluLaomAmwSd9xsPOVFvM10C46qDANYUpzycnVkNmyDNvK3dGWto0w/6jNNTsnfc/7V
hxHcnT04+rDBLqi4ez+EYXIW84z9FYmYztV+3rLXy+2niWt/YA3Nn7bnYrQM/oWqSLDJhrVWgABq
Jo+96DQ2JMi9gIEKKi5P22O0OSDY/DkHLBak7eLrQ5WLhCPVCnCYNJWHzKb7LnZNu4MJNuhmC+gU
i7s/MU/0gMuFKnOl8DHs43P8nA6Jy4k5GzZQKIwc4aVElA2ILzWhLQRC7PhDqCqkW0q5vAo2UR7A
PWSL8rU9/yrGNDiQYlViTL70qQ6LhoSlt+/B/qYiLSS6rG85QKhV5sikCxxILhziZFp0xtm4oD4w
sveEFBQjido3jSf/cH8CC+WMhpXbhFWeux+vZwroPT60fyF4RW4uMypzcseoT/AJRTtU3kbk6oCL
+Q4mtZYOieA36q6o4Ffz8u/IXbp2K7VHRvts/xYOgirCu6ciR0AxA7D2lHT3Ef5Xw+P8j/d2+cKo
HlgUl/RO5BsnaLobApauhO2j0arHNjw8xSB2egKjoANJ9eEO6ZtAvyO80TwgmRKhZdqFACbyCU+a
HJmglQY8MHHLjuzVQcsYXPrTwv4K9390FLDBPgzR4xP/zfAsWXbdKklqD1N6u+7w+kemzRLw8ilF
1jL6xjVrVqnSsnY68xP6xOvz7Gc4PdZU4O1CHBK8MO6Vbdg70HQ/LzZYCuCnFba4rCwSF1CrpGoi
U4+lJevdIV/+lVg7EuBOKaZco3sazrx1TN3K9+yL1irStwbMOXkrzhsSt0jjTWe0Zyyh4WhcjxEX
0CbpkQPKDucAvbnhqHhrZDrMSQDCp2FehjfP+iIWKsC5Q3RPkAbQu5B3p5ZyW6kDLXSEJf5DXH49
uIiD/IbJ6Oe8i/QgamoW6uqJHbZsnH5MLTbtDQlYIwQrdwj1nTFjk3YnZ8D805kkxx0ig/WsjFJe
nqpgT8xEfabdLE7kEj7hXul4wVyVuSTfjzQQ/JDTxUtLx1TxC9k2UhWPqCfLJQxAWdEvRlfaYj2c
EKhtS/EsYlsO1N+pjGK4qgDnMvX+09oOwb4IMsletV+PRW7ApSA1++sN/M2xcebDzcB6qoIRnywM
9znuGoDnhb5a47zGz76G0IRl4QFNoS9B0AWOXcNnnrpOujfChgHIZmtu9SRWAQQI75iNY1gpmcM2
X7qj1llw/6nAvzPhuiu6yi9VvzTitK2mZCRgjnsRpb2O8d6ErhGuUkssN5ZRIcQ/6P/muRb4uSkg
bdFIlrZt93TOo/QRvC0uRql+hwfq//noPudsEzGUt90+XmT1cdXVcgRnB7KOzhHdq+aUaRts0yVZ
1gOYr0PY5FTjiomDu2SYsJtebBbCWEy09rk3mCUzsEPxRbA9NrLAxB1zUbc+U5YEV/selnJWQ+cA
YCLjDtcLL1gLCXD28jqOQKE+090XsUkPs9U4WwnhglLTO+uFw1B9Ja5AsaYozeRtHditXEIJBPNg
hWwPWsd7O6nxUDtFeD0jEGQHmeZlv3xgm5TzL7qLbR4i3xP//7qNGINx/LbzsEHbnJySnxSZhOy1
9xteUPQANQccgI2//SG9aDkTbEPqFBe1TfD1iYjlF7SuvjpQmNCt4vRv2ujKq381FWkNxh3yU28W
K1gE3S3xsUGPbbXNoM82P3urTzF6bm0xbulP0jd33yGso6a7MT4Fth7PHFF2oh0oEgMipVE4VvmT
DbCFbpy5v5VoUQApbZ+Qqza288aqMF7iDKsj1vB8ZIDpEFJPbtsas3cNLtLtca2h5M89/JLnYb/B
xvvVldE23+7PGVcaAJBDMd5wRFa7CvdlMv7nh4DCHrsspm9JGtES5mryHq6qLLXDXXRHH/v34UeD
ORu2iggwRmiQ3oce7AMwL8l1Nu3bO08EAcVJfHTYZLoB0X3ok9jLuh7Z15j+6m+33z7kxU8KR7jb
IsLwRVvUr9H8vVVD8KvR/B29j7iElLC+yWfTqvQW2X5gBPt8awH8btxIaqT+unXUQ5k9C0q58WzU
ph7MUILvR0gAHzGGWDu/QF8D3P7KoYutxtOgLBK8FmEKzlczek7Ls4WfWZDlCdTUmG8MLc0joxzf
Kl4bjPeiPi3agZ1I0WfIxUQwM1wxxWiffd6s290un1Ny79uFjagz75LEL+IWO//BZ1JbSrDRcrR6
nR57dRpFiiUrghKL8dz30OUgoNXSEC6exI7YX4ecIqB5/srTgd2XvdZGvueM15R/bsdQsIixBYRF
1GnYc+ZoplJLlVAppssYTJmSFZxxyiMcj37ZwI/EI44CgRnZr1bTyBdpcDDGNFdpJQVnrSBEcdDU
gl6buSKwoBXXLSPILIvDdgPpAOPjfHS423KxPaa/qWLyuHM4IPS8FuD6iAzpDPHc3CeOMkAuEvmm
Nzhw44xHT10hJxxyearNgBxze28JW64nwh+4Pz7VvomW0qxOHVTe+oHtFYCc8tapTiUlHj7ohtbY
qP9LC1CsD0+RvpARuPLCKDtY2iHtON5WtCwgU9twLeI2dtmcftWhN+yGtFMtbMozliYNG85UFxyI
iXU/8pctwH+QRL0j0qlGPHigw211KlrzQeYuIpupxT+pjvAPVJcP73wo9jTGVpQpgx/FlfrPwQdu
SVvJelzUsWT0EmY7OyZ0tgJmgkO/BWX/XNeDGkEOGZoyHjozDwbX1Q+3QyqIg4yR754AyTsqUZjr
666WUkjheE9bXTU5KSS7MDlFsYPyhXb2cKSmhZH2SYS1fyiQjSeaeGWNMjcdfMS1DE2DdsnqgZJ/
436ZOccKTxSmOvVmX3OE/nYcCkByGDWh0cO0AETry35qVmjC55dBS5T8Ln6R6VFeOBll7jAHhQRR
AChe/zPInS02cwdBJl/NfxMIDU6yRzvkkJUmoBDy5aP3qEfGLpuAr0vdZu/uhC8yuggC/EQVrdmV
C5HcEBs7C8bYhu54hEJ+wLfw/Xpuo14Wwcc/KKljvFhF3qROx6jgHn6njqZgvMUXdMP3kGZaE8S6
8eSqvK/f8Px445FZ4GhyPDn4IboDN3q3x0k7wgOPanPBSoVo0IcRyB8Oc97+bv+t26HXGUeF1ijF
FYtbpZWUZt5nfYuQf8UXTvaw8C+hPmWn7JHcdAqptVJ2j6//xdK1cMzLck0JxPSAeqOU8GrYeeck
e8Z+K6l+FkdAL6lG2o1dGQADBWhGjJF+U0WPmTwnGPHMMCvIyIl3/3N59c8Bbtll0g832sjbR+m3
qqAHmMsefg+sv1md+RQZRoDiHMf2eZLFZLEVv5fq3QEQTgMh8qYAACJZaKFN+xNA0fLGtCT5fI7o
AfHAUyWxPu1jDptK0LYb9q3Vdlxu6FePpNTIPHPpXKg8NVG+LXXjx57nca6Nfks2I4UjN3QkciBw
PvtlC5XePZ1xRh89j8xVTcP+kvK2UU66AW5gopwFE9cYPxkPVQnHP9sPDnuEcUPYWRudaNtg2j55
9qv+o/sMsYcbKuXFtxocy1mmDDt+4MWng2tDvP4e6n3FtiWLyMR1jxe7mOkLCOkKfBLVGSsVRAT7
5v1rZbi6pM5zCCl3JsQUPoTrEcvw1te/s8OUEWPDKu7dI6Nc1uUQN3rfQCanoJy3csB3hQzKHBiF
fVr9sHA6B4nUW5nmosMuhSHc2GUzel+DJftCacKBMutwVsZJN9bWGyJqmOAKpYcXjPpvHkKSc+hy
4ANnxZjD+WNGCvliY0z6Kh0jTH+XCIZlmvsRXkkF/5sv2WYmrI4b0XdIisFuR3hXJK2sG8SJdQj2
ma2UCzJpxZNrdiPY5g+Qwfrpmj93eSp3Wxh1AxB8uv8fpIqN1TXnsHiyNZTYZu3VO0uSupfp/N16
xclSdDvfwZFI8olW/25MSOtZdX1YpptFlQgEqblGqvMU5+bv4stZnNlJshv+V3b9DWZPWYCCuaGu
BTIHwtOEv/oPDHszgvlKauj+mg9B/rZAzXX3NyKIUJ50eJ4e05yZYoFdHW3H5akCQw1lWY/kwnY+
ki0Z0JtWAIM4zf+qUUfiFIK/sETJxNqKipJm7Nqr4dTNYP1CBVdZthp3GoKjPnh2FpcG389Q1nDx
wWeH81/WtBmbdutXNz+ZEzO4gqpAW7VpBXIoYeDD2ryXsUzBkf4s+jRhbgtmEv4NIiIt2z17puyX
97ORtriltPVZzjbbPGnztnffbhCIgqhcYpM7gdcZSbn/mf8iD1wbMSMn3oJeztr0HRKpLVXQfr4w
NfsS1jEBXtiemIC1SFP8TeMKQOGiHYAQVyVuNxFWjr5Y7PnET6a454VSuLzfc2sjNDM/e67abhxj
QbMT+ToMb4epQNuplWRIQ8j7goOLF14OCyfBDd14Z94WxI0WbEBgEbpEboTHG39/mu1FIMPV1yxE
UAVeqZQBTcCo14AdZt1FcCMqSOIB1LhFUyZfMnAwvjFtQ2hunGgJLm3P7l8FHzafwQwKzsZGWuqN
qCSGmwvFWaR/K9U+/ddhAK+jleMqhnCAj/Fw60aUr4GtjRinTYgTlWay41aBqKqDrUKU8RMgflmA
cTTFCtfGIoU5sHpMZiSb+/zGPRHE3iCnZOa4d4ZfW1vM9FbjVYbj3fUV3lZvWnECfTAOqkvx9vRU
M4/zKs263I2Rx+B3/uFCqKrLgcWpvwSZ7h965hhDkV+Rqxd6S27bOWjiRypndwTyDxS9tbW4bVga
87FA5mmxELIfpN69K7IsUhB1ZUsQ1RF4dVTubfrlsne+US82qLy9KN15YLLAydLn/aTtRAYkhj/O
/kG7ss5vQeeadFo42e42KfQAnsKUkhXrkk2HFoG86f2JkzrZ69nEAz/+JoJJQP36cJdEiFJ/emVX
AL3vTCPYZipB30mByI6h5zuzQx7iXOlsxTzNiWZjO4jiI8y117U6W7n7KWEp/7/qiD3Z1r+NFy1N
/EmNlkQ3RsRfGzMR7EHEFQhDcpwgz1+vZTTih0EKXdq4J1yMwbHg7tFdNltM3w4NkOlmPUucMzUw
zfvksTrS/SFCLuUeQDP0dY0E792zgP/pXQCtCWiqQlBJGILRkr8b8nyeAqB+aK0xojWN5rHSVv3t
GwftGjr0y96F7rKNzWwydQLvJRd+lnE/LdCywIz9OkaaMjjTDZUJo6COJc98+7jXMMldX+U7bgSh
cK2QCM+LrPuFJbd2Ds616HbGv+nF7EpEgwy8L5y1ohh8qAsQWr5ssZl1a6gSpUyTKLoo9MPpry8V
eEDyyG8eBn2rPJLHRnkpzV0sP8f62r2YxTzfR4PW5e4Yl/ejT0Dr6N2FDglVMsOyR+FcCRr0gaq2
SSL6SfCq5MR+NRjVb4oxeGiXI4qK2daDcNmG1jDgm9+ndPhiXG69JgUFI1EOFQzP5M2hAKmgsBR7
OVLQK5q+dxw2HMmOZJkKYj9p5zl/rsVU6Lgyf0Sw3mSk4BgOHhNQo8dlWJEcTEKy4Q6bOg5yzDfj
T4hUWAHDKQ+a2o76egNnzkcVJ1lEaDtKGVBpADTZnAJcVgJfrafPH4bRtdd6ufIzQgWYeegEjHVU
0BuMVlNKPryvM/Y16gDnBrBUfBk1vuJmU/lZAhqbsDLjw/H+dQbfuaoGPVUhCSdky97ds5EsUNGm
5QdJDRSRbuONkSsox+FQ2PvyJX4zqc0xLEHYxVXVhFXJzWbThHLmIm541mY9lKUV+GcELyu4ojW8
m/Ffbv8J4u6y3xJ4uYRWCIkRq6NhVuBM9S4WRCNxAyh8oX6AuLzj8NzehVQ5RsCmc6YyaDUxEsW6
H5Bj/IlIt/PW4oRs5CrwhyULNMh6UxS7TOPlvRUaEVqfj8x7xkh4HtHRTXeckGvOIlGNRa/YhXgB
zEJMcCuuiZr6g3Ny2OAnQxCsYtLb8qxoQ3yWIf+sf0Wde3zodbw8OzQz1dOPEgQzLT6q1vbKUp6d
V6dbMvsITi1VxyE2S8svbb7yH01ETk33RnlLPUP35X7usFVytlGOroXYRJdZScfqW2fUF+rSejME
ulNBoAwrlUQVZssvCywBQmSBzjVqTKifhMvaAkY6UFuMmw7RNX5XFEBVB/mST2ixS13FBkwGR3DL
RKf72i6QvkNSg1vVFTV5sKaB+474febpj3UxoHKRlcIxn4llg7P3dTOR6pbgJL9s8h84RzFq+/5Z
xCYnKt5LVYBe0VFlx+rVGcj5GyQCtLxoXFBMN4oXsn2Hp9r4G4VxF3a4il6xtlVPFvIyX9w1BXm7
yQn8kNuwciIm+1sUexQof8Gu18jU8m6cl00sxy3/C6Eo/185clqTMGa58EgdmAA2RNAGHEanerX4
6LNnIXh9yhKanPBLAXEtjMcVLpKm97AuDVi7WO0Ey2nUIOrWjYr+5v6iCjMqXZP2ipP6J4lTPXDL
vAraarO6Yqd/SXVfm23skI+9BOVejspyJHpEAzSkBktGwMp7sOpBbJMEA+B0XoJTZjmBun1AWZLu
ppqoy9Ki+UVFQwmHwdJhp/f5ZNmYkC8nGPmZEoORRKXZQHvcOmXSWMMVeTVKEjbcsqPJZbM3d0+z
gPwLgVJV5i3c6+irHJ3nc/zCiX0ttHPygRS0HXIKnHwT9akPIJWkBpF+QWz8dQRFibriUS+Jafm2
BmLDvfR55sSElqU9pQbY2tRv2Mvm6FFc/C7DArtgtgQPyuqglCA73GS9p2TB39Rq33j0Fq/as2Rk
GejwXtdcQXwFuFl4+0Qm4QOLtLOY2UHes/iTtLuQSyUnhcBj+LZYqy8tjCHvPp9MKdsdLbelvWKW
mdBcmkd+VMfbTpHEMw+/r3Ui4ztyvqeSBZzSlX8k+bPtGm3VinBALKKI9ckFcOvu5w3/FIuwrasx
5gjI2njx7AHxadKybbJJGuPQofjHiBccmi2zaHIgImbRU1GVG/ME8WftaElzR3gEoTBfVcJQaJ8+
SZBrU0LUl9PCaSHyF9xrVkW6EZm6i4OqKlvNQEVE0lBqW3/1c0G+jw0PzH0WyCoe8YT/R1CDScM0
owT2h/8+fNRf4Njs4wHIlgTw8KUdWIhZsu6roTy8iTReB5+6DmoNIISdvv4vW2Kru6Qm2zvFBmTf
IwiO7R+ZwD/4h9ka5lmCTMaAYuizhuWAjsxVxQ8wpwvkFEFpNNxyY5ppTLKQdnsZRy9wewrFvf5C
PToLSh4RzotGluxT3rYfby9/szowvlmC4Kh3b3r7kBiMQ/f1Bzm5BU85Yhlz3LaKBd0FTvofxn/t
cFe6wFq7raJESu+6NXN9vwRYD5YKTB/I9XDvq7xsFN+kMfh/8ROspjNkKZQj6WIAqvpDDvPYcjPT
ekyezJmSWL28R5/L4lhtQFrk6NlMDb1N127qind/N5IsZoP83lK87RJWHbLCysdytpVvCz3WtCim
CFMWUPGGJxNCeDlHnIHOaZGyLCCbI7+wzJiL2iAm/yX5eXBc4TsXnDax/Csx/X0N6AB1In7JZb6T
zxhy1v5v8ez53Jw8XaPvDQMdgGERrRj21luJYviaDTqF7Q/FlJ0mSGOkPVTZm4cGYO+O22vJlvNp
vS1aignQDi4yPrC7aPgW8vYaGE9XB/TP6XuXTLCBp3YPo3pKtkkf1s3hviW0DwKAwyWTJ8z6SlGF
+CJDJsi9N1vLsz/JJGnUcThf3KFCM4cvF6JqAmzCOuuSZDmljKVuIz7NNKi0/b686jekXXNMQ86k
7O1SMhz8VyM2XT33TCEkn77s0vqRbLiq8YlUvqcNXBow8WLOZzHeORPM99rmmX7DLNBxzJnSrfKL
8YSXcqgF5WhXgcl2K3LreGqBldeGG5tuBnLuamk6ZxNuYzZZS08ep2Ayxj2iYIrO8lVzrkfc0/Ti
WWvg5a5f9fscV+Bjre9Uj6mygApWt6TivCC3PPh0hYKRdDairi28/5A5ZBFXkEAM848pO29tjK2u
rPtAcC0x6/n0jjGXs6XBXeTYZIQ/C2qn6WxPRE8hrro0HYXDKqherk3ucodpcoQ+V42CkQFd6QzI
PdMLyjLcwDm2JbZSHOvUSYbMs/s78S+IWyCtynw6EkCEoZMRk9KrfexEeQUUc90MSvULHnQHLJEo
bM6s4NlrlfbqpHOu9FtliqpJLDO88cvcXCXsKFxpYG9GN5McWq1e7ibkQf/Qc64Vg/XgGrEVSXq+
5p9t18gz0mpM9gYfmk0vm9nmk9pGh1UC4xbiVOLRkE3knfDOFZAKoOm9g0LRqReIvy07QQyuIc0s
UM1F56MqsvSoKuCoA3ZK6eRmFppFQYiJV+2vE9R92Q7bemSSGr/B9xIeWTmfy4NmCk7Q6P08RblW
rLElB9Af5hB9YCHgz3b8Ze3UxXT1/Ha5p56E6f9k77H/OBe+kSqEmiG+GX3GV+V2kIIC1k1+aHuW
7SiuxU4+VyPT6FCk2yZK46X3oPXRoOvp0K46LFtwWsNgqxSDfi0ZG/Oztx86QZIYenwKBKzFywbi
ja68m0w5LJYfiXuJdh0m1a77xwPhCjnw2kFelvqbF1HRQ8LF8iRCCsb7sfPjy00F63toRsszxH4b
WMvzXmRd2DjB6cH1AUKaN8Jk/MxuCj5/ZH4lDGFtYw6oCTQqMBR7j+WS0sFKC/J6/j74XZXOI15O
sZYwgnKMR9HVHLC90StWsj0QPasU0L0cyrT2eCd7F16e1Qi+g/pdyWOP0dLo7010TL1Jn+Ou8Bwu
w0W38N7sYtcfYqjq0Ujwa/pqtWbdVqgJYueIpur6/cNpwDAO3xT5nme/DUjy8oz/9Dt9SW3reb2j
GiSn3rG780kcY9UQ1XWG6mehI0pkf2EEpUo42whzGGhYUJElOg1xatlJd3rSChF30E9CPa8poRfn
oNbtfzJclHoFcuWwnvQz1rUBnZ2ssBTsStIBBWzaXZsCsxCFyfzgVL/mOPMnhqBe4nFZ8Kycky3X
PoiJb9m3axhtxHJ7nxt6K50Zd/1XSCF2pPd+eUONj+B+Fba4nmNTlvb6/G/07znZHgmrFaQGthw4
CoDVXnXQry6YrI/UELWkU4OEbdRrWFKs+Q5qybmo33PpX2ZmXbTY6iHcSMKyyrEGhxKRocTPeoGH
mkZu1O+XI+ruOU+SDR1L1RtZjKClz5w1Ttd/1CI0+S1GWETp6ynB2ojeE8JXwLmpP4FDc9/3o0Gd
NRJUi2BPTkE9vBOMsl7FCD25zx3y95censIuUOba612zRToyV0e8ApRsBfA5rBFku0g7ElJ4Pccy
n4p0ahQZXFdIV9pnTfiGc0cqPt4CtAqw+tiRiAEv+Cu8DC8JtCbosFrQL0WH41F+Ohzoxzke7Fpw
RmPVQp2BBP3p2Od36p053OC0K2Jkbdk0pJCLt9mc2GEwIvfrUb7llMk0DVOx6kPQCHL5BbgfmxrX
nCVId71z6fTqblDq5iwnEZnCKJUNeLxJ62BZgSsOeWvgBFQf2TZ2qL1IqPgWhKZV9P6Ow+/jIdV5
6QKdWcPQ8oPe3aEOULDUVNfh6ojEOt2zBOV+ldxK0SIp/58iDm3fzOHrGQaxzKh1fG1O1CuYQXMD
b6DLfKj/QaNjF8wdnOt7ni9rwmyyoOObWXfMi63n7486S+3hX87WnOLZpja1xkae21V7C7XQ6xRt
wYLjWxeq50ejA9hIJRZ06RIkxEcU7lDABUaB3gKaCzdM32KOIuFGcMh4ZNMgeR/rLCsQ+0DvqN19
av637K7PwME3SnqN17c8bYZoUEJPCDl1JrTdtDYzA3OXL6FMGVjrkYnXBm+VdMt2J1S3PoTVXcN8
MiItF11SmairYQ1v744LmagXMP57Yd8FnhFBhCuqU4NQfcFyXBlW+JdAJwDYErvTfij4QtUoU5+X
EAdoPJ8tKE2DSQqEMWAfpa0YUYP/OsTdC+J8YE236ayFy1BMRJm5TMaNiaR2jAIS6eZKm2lg+A0C
PBfBoufsdG6INZxAsbhUEaLq0owf6V1VZdqgOeS3iTkrRuG+OChrMLDCwq6xZwK6oFIJe/kG+yzF
7XXHEhIEI3mOkwd1BrNMiP3WYyOp4a2iAFodVhU1ArkHVdyFVq5MVLAsQ1Qghj8o5QIgEcZCAQ4w
Mi7x/L8VvqZ3vaJx7pBd25oGmHlm5bZtOG/xBgt3Iz9UcCndHFahu5qVppfob/ihRm7Lvc27Jt/e
0EC5auqU+ErSosGm9kTblo5zlgf+gs8ecrFl9PqTKVdF2SJw6BNMgD9wttBlC15JSYFAKuJQiI4M
zHEX7/VlS5MHEeavdSbME21kFasAlOI8TzpfMCXOqU7HvbWi6lLobOkl46CKHjSd9YkXi99Irbx2
Eda4Wbz4yfMom/OYBz4ITDtA/w5x5Ad1JTgAzS5cCVKtDGPtvSs/IkN4/9n7yCmypgd6W2GXUVcm
AqlJ/Pv9y8Fqg6o+VnuzZLXlSp+Qd4kQnofk9mDkq0GiSeWO4jOs/Ggh6T4V/p/wKudr6e+zPPuT
JCt/Nk6j+4KoLVaNkfz3f96/HO+DBylsXpQ06li1J6+YMG22JybtaeQbpkKULsC1WY1vXWcvKSok
S77nlV2p7q4/wxGqHi4sFtFHTL/YiiHRUfHj2GGo0r1f5QZR4vVHPeBYhRn+gREd0Usb4RSKeGSn
eDKqo8Jqd+heGeF8yMv1z7vBUj/LKUCFn0KH7Wm4l+kQV9UhnGrGsVzE7rr27XkVbIXZnB31cBsf
JakqfWonSA8xVnhYNUqnI1WaVdfGYEg5OWw0Wjf1Ixs8IWt6eE/YpLsXV+7Sg6a7PPAqin0Zg1AU
mv37stIbELKZblv2p5yqUhGqLP5xsg1BvxVdLWjQntDM4va3NTwW8zYFrKly6orybdhEve7hapZs
rebLdbeFgL+A9bZj4Kke7awkmtHNSLwsE14bbgs2iy8Ozm3dCeklBFFE1s8MA67yAj0Dus0FtiPa
RBjZO4MzgrbpvIBLy3Hn5gicJUZ2ArYMxWbBii5PB61LhZYVAn0k7r6a9BBHhOPuCSraJ14qShzZ
AI1olvjJF4rIlC/dlJW0+vIXqzuMRxZi9tDBdqwXTe6p2VlTeBnQWxXVLvdZgDpRBUGZnvfFCiAg
l6dSxw0BWjxVRLR6RQiz6d4lzUt68k70tz61GhxIzSVwynO/Puue5/DKFynYlVteyVp38/wv/e+F
+/cCLDS0yPvkmAJZnmiln/dlImsvpZJqpegaMnQnP/vn27aXn45f1VnIdhXNYPf6QqktY10pVDY4
wvOT4Zn/4FY5CuJTPBHbUOZ+jSe0OxTbh1rQyyhAzg9e+r7TShHUMP/oGpgx9iQYZq0RnzNlq8cJ
aaLy+T6XXeHqJhr4hGQ8qB41YjPA7w8D4hdji7u78xmdiLGKC9rX104WQbbRaW/PeGL9M65A2dK8
G7KD5hgIWZzGo2dM/USYe9J3fTvjN11pbNJ/5xLo2vX/3YqYmXIgtI7JO/OBxaKyec63yDb2b3Mn
oNquOwJJEq+jktBrI/JIvtwg3/Mjc0Zkb5NxlcrUP7+kEv0k2DsGxPE8TBkmuSu/Kq2+vpVIzs+u
Pvab6KVRsj7qOgQmFs6irMmLMaNLov91+hO5tdJvekNsE1+x+euriSZDcJyj7/X+r6PxkjV1+MiL
1gIiHXv4K+bOby0KP9CfhVyxR09gIKr6zpNTYXVpWUNafCi+N/A1jP0TdDWJw7Cjt9SAMOiGA1zx
rX9bQq6Gm90Pt9E6iZRP6beOQl6RY74Mm5zj6lTqll7p6vp4ZarqDIvcs/Hux/QY0YspaOecz4qh
jtSkoYIWZ9gzz6TT3LjBrzT3y8tyuF5+eRzfV7p1DbcHfOKcEgLbmjlHhUNUoGYQdGbpjVhLD+GP
hnonkEktVo+GNKWernAah24h+a7GV+GxIHRUk7IcI7Wuk0C8Zf8EspyVYf2IHR2CyXhKxE0441Fc
Awx7fwQNXk3CA+CPjd7Ej7uQTqvpOy3wuQJKggeC9xpiItTK1UXlJxiyZDe91RhFN1vyOOtxnvJz
g3SuVnp1j/KMrDSg2gpyYG49VPsV25YlbHTNskhRDn42jA6ZvQ4UmXZLUlYTe8Uqav9b2hMwsPmQ
XWJ76tKGu8YjgG7rdION3qJgbswgctj8cC+6lOmvBzRJsZGwPdXj7mDHRmFZRHw7WdQFKrcZaWZk
xOlZE7Q1e2qMse8crTt8crDSHOfh7Oa4GHelAT39FB2xflbYlNTyP7VMNNXb3zOa/SGP+X+hBhDZ
AAJ2kFSwGgQ1qck13mL2X6WMOfVIQVp4c5Nm5ru/PY/CgaTkv2wphfTBxwhh5kCSSVJrb7tN2t1a
Zn6BcrJN9IIfHqafAVotpXKtbs+L7RctlvfNawcBUAU3x/AZPSCRUPc/jbGEv3EOwK2OV7/T6DC8
7mnVZLUx24a2BWeArVmcbSPNaOyliKiXiHQBP5O5wkC3Akiz17ZLTlcGf4ibdoP/HZc2oA5DfEf/
G5OoaZLjQuFZTQ935bpoBcUEWGiRCHwmn+gZyaydbUzUvNhaPrmPhC9Qy7inddVW6h7RjMAbn/dl
SsFdyhGw2Gco26sSFMpWuy+c7Jf6qwMuExfJmAK9i0qF+ulGjWH9m1/0RYRP6lmpJ75tg4PDzHlC
SPL/t0rlQPyvLxm0GbxMFc4qafat7xoT7ZllM0kmy8kmFKCETkchQXFL4H9UNsb7MRC4iihuDNuk
JXMG+7M8FK2j9HgrAXfnPiy4zBpNeQOHekh0bup4j/WEX3u9b0mHMTxcw3fAfkejmGBgXG1wJo3C
fY57e6PYArggsrqIMA6B2Xb/ElSQZlEPEgLJlDZCv8O+k6IeuOlsSnq2p80VkuOLEDmIlctB8uS4
uXD+Yx+VSUOBdbM2Oxl4uB/BO6mONPnCeXIJJhpmMo1OqB0qlbWfLUrUv8q8qXWO2s/gGTPd+pCH
Aw3mZ6tDJLYlkAk6FENNZ4XAViZDaFqQrvAPOcCm3/LOY6AwHJlq1cwpRlz7uR+/ALW1mDtQSejF
KrFExKJdl7Nh72HZh8sayKixTArpKgLbEjlWpRzQBBY3yw331m8edjM3kasG9U9+8VBBg7d6I0Ob
jBRU6XC2ZOPFJ0asE14PhVVgNKZ/rN1my79102MF+aF3aFczaqA6u44EzVuyMVyKNgUA/ee4unHm
yei/Xr6O23hXvXlnTBcBqh9oAeWp5Yqviv1CEMo/H01NhPW63hemCOWV9SiKqICCZ/D0DwUBoeVD
8iqQKlI2KeOINLEItsYEs3nxXu1iQWrsgxwblDvFDKS0ARBfa8oVwsGpuMIGjdir7ZGDQOpprnGX
fu9GzPIhA0HeQLW3Swc+AnalxQnUrrqpL3vis8V8GH8fsE497R6KqLNJS7xTC6X8URAmCE0+hTJr
+YqX/HxrCA9VNkPDBJRhc9SmYSSK2tDtMTpBkfVsGq9Q5HiAqkN1m7ISSSRtqARCni5sf29RDUEN
j6pv0QHxvxupyuoO2c9o89RX3yCd9504cKRXVP6HrCNWfdI1R8t+IgNmf7OatKs4Y1YU3VI5SUxG
o6NETavPfjq5IjkbhDXta6HvirOOgbw83/xfWFNWN4lBofD5RPdwfXjfUWtyiY/RywKr6SgkQ38k
mT2nzJAiYkJ8xm87hbIrcOUrNuthr0NiXS4DpuxoLb/iVFnlxCVm3yy2hCpk9oY7OFAZaGKxunSW
COTfCsWP1Qb8FtnuLNC3ogYdYl68YYkpVDzVI4gglLoqlm3k1/CQP0aZtnTtTU8ax8LOBFPthTNM
U+1zH3CiFJzZw+sN+XlqYGXL9ZiVmlttaf1mk4bgGZivZ78RpedQ/jGm0B7npcm9wZsNV9IHf+d4
uP8QRY7Shse5v/SjxFUNjCW0hVfNFzsqWftSmuMBjLHYpYq0x6cb4pdHAiB3hoMWeGgGatDXRBpm
I1zshPCexyauHm9lEDAawp0MAlucoPhu4SEAO/MoJR4mVe8bmktoelih3AnmhCS7COKDWYkDHgJJ
/yaHykETbYxarIgOgHjfVFyUuLLp24VZge2QEOTofbz44e2xvAgyAk3liqNyTFFpl9PBJ3ZKbpq1
EOJIEqbwZ+LXYCXqXQqL/v4qRnBZ9Ofy7XkU+eL5FBYPeAg11SjYtvLVAMxh5cIlyd0JpAW79mGu
jdDSW5lJKxHPiXBB5ib9PVa0xVc0gPFFx5xytsOiIiJ4Se2bv60W+k6OuquLOjsctZwMN/JqnZ4X
mMcqrVfK7U0LL1HCNP6M7ak/8A/pQRH70PDCJJKBlLCiwXosNwv/wPY/gU4GbZI0YVGzrHOO4YGt
nqkcQ8FG82N/liLQwSQgOHsLkk7gw8yM0gEqvwO97NmvNGTGpWjKLScZzLqTH2/ek0u1BRnwZopZ
mpoeGMqUZ+sZXjzJf+fKUNCh0zege8Ypxp0JgEsQuikAH/uRjpFlKVF8//sY3UEjZ4XHEqgt9pwU
4eIE0Ntr5xpPSvh6D3W25db2QFPHaHDRHh6olRH8IgZleuZQCbjtKdY8xQF8IbLdA/a+UvItMxVF
hg59+MME9DDaTOtOOZ3WnswSIkNQQEZv6VjZwWtlzpnOPR76XvDMclgBGpyIDv4v2YDKbj9rtDaN
ONXKN1tDIHOtgr0gz4wf7L9BRYeG5QPJak8CsH7lgnErvcO9CSKP9W7cd0nF65+Vjdcn0l+T7JF+
cJ7vOrD+p5jJQqVyQbI5QnuVZ3AEU0JYoHfvM++A6IMh4k20sLZB521n6WcxH4279hCZeTUJJ7gm
zRYw+uS6bQugMI3mpH9SN4zJy4ve2Wd9vvBAwbwiBamscDeLQneRzC9kLGFxdgXV8ZvQicG7qDvk
CaoBfaTjmKhPNU80bwW6dU9lY44xEQBTP1hggoWFbN5tVEsoXl9r0Ke6cZA6E8HuLnDEqTFBN9vw
0CYPSRFvH7rRW2iBUHzs/+/YzzFyF8AVOBiFNjLDP+xXWhDbzVi/p3z26mrCihyDpOUvXeQkye14
BqYnOYunQHnFaql8f+FcelsrF1e6Ek3eKOg1/1iAJPr8XVFIAc0dpCZxhwKPJBNt0iMy4E2GMD3R
yYkRN82aEJWExDbCgzJCWGmz8bYhxQPXZAnDdKW+dod/yT6i1NkQkgCsR08JQvzGSR15KRhwmDly
9OlJV+5nTk2qNow7M3op1oEaa/OIkgXyUwlX9Ovj3wrloyPVOK03GT9ClDnl4Z2gmvDUjrxfEz7Z
LHHSuOBJAhGNnXiglFIG5OikWrQpvKgVbIK+B2Uzfm22fmH1I8XOybAW+SdaG2yitZ0C5WLQ7bxI
+KhWwl8gNZFnV7cLiNyc5wbXWDgZUHUIJN+vWtg8xKNy66EtgBb/bhJzlpHxXQCKPAFUsmNlkLHb
baUHu5jIkxsPoAf3eEfZw+m0m3IAvGngCcn5LtHrpuar+L1jo8L6L4gl/DC0zZ0AYwJ14iC1M/B8
w9o6tlm1lJ8UEmbiuX5fNJwoeUbNRPTuzKZMXdaHWw0VG+lp0Roo/lnip772q1AtnV0ncYN+h/qg
92CyZ4UH0R1CSuB+LRHL5885LGiZbQS13cVRNJlVf/eSwnn0CCJx8l94OgGMXRqzRcPAy5pL5H0X
2i3mTUXCaxhPRPjN8/pO1vB1bn4C9upF8/8FtClQ8vIRA0Y3VXovU8a+ys4w/qySz81PNnorFdL4
XV9XyEdg/eWGA4ogJ5hSyQm4XX5x/F/zF4ABdrkjt94xE+25WPxyS2j2CUXt00Q/Y0w4fovGHZrw
xIpHur4DoM1/I1lyolyJ75k64KVlxu75wmxkbHOK1Jr5jSb5MTBRUMs81LAdwhW/6HLjYzffd3M2
sE3mBOROrf75kZiz3t2xpLs0aafDI8FKePWgggZNCKe3W+w4x8i4o1Fwb4UyfHDVyvxF+h4UUbIX
l8TpZoCawvARhNUaIX4OLd/OKKo95tHh/UWVODOqAOxEwL+grxNOE6xYIaQZO73uYFKhYHF6wBNN
ZqR3jD4+HKdHCJ0TxPBDnVBPVy59EsmeHJGU5FQsavSNGUml/GJmF8Sp9KXZAe79+Gju40L+VLNb
ChjdhKhxQeDZhnc+jyt3EwRLdOC6v/jA9Xh8JuZDDU7DUXj6vt+UXR9/CpEWHybMkW6Jgln58wKA
Tzyds+3ZWK5OLv9gCElRarq9HT/ZGaBzTngumNbwmdkCJjAhDWh1K/z1EbLRAzdtlWv8sRcH/r34
OM3j6d5m2goR6tv5H+SHiZhyusbDDCEf98czQp+ssZDMnEGxp/u+OcaKFtqzSfQm77TkLCJ72Nn7
og7KMzV6c0q8Cye5kbO3bguZ8m5l027qzLfOP5BXs4/Lbr6rveZ9XkGS2VByuRtgFbvI2Z1fBf2r
3mxCsNA1tnsI6x8NKDPalP3AZUqHSG5Js1NBkiinb+XvlSA4KxMJLZ6y2T9mXl4JggKoFg6itcJz
/bEvo7hYFQZA7aEYoUY5dKZdB5n9V9O/GPb/sjg8QXJC9ecR7MKEo1awyqNroOgEGDfLYDF63Tqn
HWagbDTyeZw02I1bezJF/R4fv9wXKNzg0fvpvCHktDfbEU3fEq81FA7hKBeYKeoUgZFl6Pj8GQpo
4l9QHUJ7zgZ3PuV+0Mu1EjBZSdg1mM97GE/N4+OJAOU/M+DLTExpI3xE3TOWn8M2oJydYAxFW7CN
0wbDH3hjnDJF+jZ+rEHGuY+TvMB7oC6RpC83NcaPDl/fQNp7xlhBkaBrrW6+tu3ikf2UE2q0o5/D
vAjG0KFvEh2Sbunv5NMBmxNc4bajLywakI418O0b1Bfcad+cfNu8r8x+3hLg2LudFdn5fyGRC63K
rFO4NNBVle+pQvHRCGNiAiVpxzTjzAOhC55BUUjnhU3n/Wow8imMU0GlNRJvaHU2RIb8tELOT+EG
IlQE6qk9aW++mkfPPEQTIuKXvN+efKAIkIHcJ+YrxCVgV+cJ/oxrEfKYJCy9BKQgKMI80iHLF0X9
0oaFI5DS5+pYAcMk7/O5L6cSp8kVovI6n3oXHiPz1b0j/e8Nq5DVdAALdU9VuLJMMnpMydKXXkuR
lVGxcWam8qztwVNJLA5a9Nzu8D0dovvckk9HVDTq57fZyRHNz4gZdVpUcYpYj7qTjNtE7BNw9RTw
hUfyNX79o19Tjye2JMNq1BU4aaP/SvnDEymduKf4lOgCz393qqNx+jw1i1rjwyYTAzKJmiept47K
p5blNJ+xYxVghnXc13RHLtGZQ3IZD22W9FbQmlHiIZFAZbWQK/j90cdnC3HX1ztzrSYh6WJHdf1d
odVCfHUXPmEaw3MbqH21G3ovC1ol7fBpFQ7bXK+UtIaXbSz0HpmjAOkIc722jadp8bYgPxUokLXE
l6eUfx/EFKTeNUqq85+db5dNOHdgEJPDc4Es7m3FUbugfYmp1ldj/evMYmEU/pdNEVnNIPG1fac6
8DIYi+oyCLeHClTa5Qywrt8RKw57e6VemFPxrjnxcaa813VLTDjSfHJZ5h4xTKZFHYWurcaC8amS
GRat0ti6CvVtVc39WnBFCYDzFGcv8PvvuBeSD+GHy9vvfs/QsdeHN1vKUIJwiIkGSHjVeSERIM1C
EmS9/+YKemopkungEiEv9235LJVcz7RMroocanhDSJ5AG3hWNh8amz+Gy/rCmlwpDQs35G4d38Jm
oB4iWgAyTxkjzEJnc27P09W9xhV/g4Y/COEIBm6cRtjtGGI1Kh7bkJzdxCaLAa5H1m689inZkIWB
nLKcThcotgmdVzBec9Rtrc3sYtiC/kDHs/ek26qiCCCcfMANrNbphiZCK190E09QKEqPckysb/Sv
v0Q3QqpImvuav+G5n3u7U0+7cJqWPoxXDxAmnSDx+nuMi6hjGARD+/v5FYnrfZGkxqAtw031QHK7
1PF8q/r/FqwFdkn0Xbxgh9opiNoVdcJvSY3N7G6vvuEL9vDjChTe+NwPcl53OyK+/shBKeq+uYHu
Nd56ad3rBf8IanP9g/w1W5goFCZmD41P0R1kgpDJAUUdrc+ekwAsSJdrzEOfCeMfUYUFEr8EFzW9
UOqF06txlmfhHoKPEt3dfROQ2Rzp8ZVvzLghGcBe9Kjd09417dYOG9GiNgwoJDfnJmurSrKAG4if
j8UBlndQtaC/FrWtXhfr5dbQYrd+0ts3fpC9yH/g3T6Uq/eN7ijtH+uhRx4b8IzkDRfTAlVd44Yu
JxLOfJF2euPi0BMhS4kPapgaz1/07H+dKXIMrGUlDLSa4JjylLZFvPW12m7TDUKuGS5c8G35DIhM
VCNV1UmphYCBEiFXy2VOkMIKuKQOUyMRv1DHNIMG/9zAIFvX1+IB1XBeRNU60p+79qvfCVc0Mw3B
n6UAMxML1i1fJ6gZLG7qoHKUXAcmWsxRCvBOim/vG+EqTABiYTepsd7BAtlOOueDPHp3lbU+06nw
WBzVwf3NjMHnQntaqZSBYOhpD+ytXgotWNd49aIW34voiJYljHTAmvoOlqAV2gsYLaQc5Dkt8GsG
wVJ+qXkoBbEiwxIcjttIYQLxlo4JBIe0qXcSpV47jl2PSaQ0lQH+AyucMsJmhyyfknkQeAoePqJC
w/Y3fPiom6kHcRGn6+2ydqpZsAWC+OlC8hXzjlKiV+xQ7VoXBbKFt+mZwaxMNYnFl5fmd6lycJN3
CI3cuDE2hENlgJB2klyAAbG1IPjAOHD+eUW3RdYfWvrxrUe4JQH38J59yPgnyfiLkkH3dTEsIqby
Rph5wq1VlldbjXJCOUsgN6INe/Z+qJQWVZrgkb/GtkxM6L4T2UMJJP+xny/lXJIu35iV4+vCQYdn
kV6DONWXUMioVE9KdKOB3YTQOd5K+y7MycYR6zBtBNWaVFISJysUHWBdoQUECOjj0+sl0S5yNALk
FT1l4TI/gAN3iF300xVTFSvYVUCiYK19ly9DcwebTDtDVVObpNCoQNhFReEB3HNY1CNxq/RLk6Q/
CxwSvPWgyfrMMLNWn4F6I2KyLtIMxT77LSbs4KbfuE9djZ+vhKUDNVQesCEgIqfLa5kor/C+U7GO
PdrWL0D/SWQ6oy7q/HcXrgPfMUYIlLELJROxl8pE60FHT++pkAMHFmJ5lGdtAervanKxlTKAmNrq
iTesQW9KUv69ti+pz/mk1FeXPU7A6ZEtb7tWDBnKRWqwfoX18wvZpW2Sv7amE3E1e6sPVakOi9mq
KuD1xpEB10HUVT+Qf//CHuKUORWtl7vhc2zzShV4H1c+FtWxBeZ83Gu5Tk9dZXcpB2Ged5PUYC58
p/mx8awjNvGTlhcdF4Tx3NkkJQ1jenkSUgslEDGgeGKDPzfa0RZM6+zIC1mDB6Z/JA8vU+6njhnp
shlyD+lPmqwUDvrTTdQXk5EKdc84/VuXzWUT+AWwJOOlsEEwC5PR+ISONMAGGl9i5ccamFNkBU+T
BX7x5fzH1tO/C6fT5fNelLLvhXffnkVm12iWh1A6rje7R292SLptZekD927ECTPk0Zn4i3e/xDPu
vubcB+7Vq/5naus7cL35OdGPO8bmVpLZkQ9F2MkBBV6/kCtfGd2s0NpSIkK0M8qLF1D9TT2DfQW+
xcP2mgXWdyImbI8LNezm5T5ZxtgwpxWk84+1Nryp37Xflrm6wVQWpTstRL0qz/juMR7Xnmh+WYh0
Lmv3U5CcWUL4YnC9CU51vjWe0g6LaJmoMYXbo2cT6OMjCpgV3JbSu6/sccOYr64Tpgu4+FLSNasy
pnCX5omJe4Fr9rSSPHR79ryZ1BtvZ4/J2FgU1TVfgd95hqcefWjLc52g7cMrJoISXT7/G7zmbyvY
tiXJQeowdnTS5fxnLlIZJyNUkYo5uLhsdjFiW3xQLGs6syCdonqPZgPM3tVRvh/2Y8qIABhM6KHu
+btI5qYFWDGXYBFTEcrMlCFOrK3KLRh+ZJR49touatNwWgeqxeOLSGaW0GlpNFCcicFpz9UvvoG0
Eu2dAvDA2PeD2yy23BvxLrlBxfRO/xNPie5Om9czL3Pc5B/YClJT3gpj6wpKzxWMGyEA1ADgGWW5
XGrBfeN3FiSWcfDyfiWQrjUgq96EpVQ7SchHUuCt1xZBit1oU1U1W11uMSigD8Y2u5+igbw7PMfX
8jHIjv2f+Ajj90i2eOoOnXF1wZZLjLMsG3TEdxHfZ1LHrPv4lvR225fYr4MjjkNPxu+BbYYQ/FLU
rDVUDLSAwxl+45lygjZE1ynpKbZ0BUcgyvmxSNdB7gMiU7kWaFteoApp/XGS3cMHdDwZsqz54P4g
XhSpc2ncZNr+VufngueI1RoeGzy4edpU1+1xv8CdaJ5d9zNWwHBemn6FTrsHDu37/YfgyEC2Omll
P/ze80ZMGdiD/1MQ6GSXtMkzmLmbVJ3qp9RJ20fFHVD5bptPMxYptBCa4MP3jqr5iYgGII1+oLG/
5CH/hXgSTbhV8Icbp3nycTy7e41THipAmEayL0aW1ztPsQOSTWLhn+vzfhVdpxb4/XRDf7mv1ssD
lhdRKLV3m6iBW/tZQn2MhtG3Ql4fUx4+JDrcHrM7ffq1sgiJnXgr1ZjZkYFr12GYvG4s3ZxHLPSI
NcqtdaliONKV+vLWd1RQ2s6nyVwMhag+Gi/qdJUoLJRsuxAN/OSaoEtkSEv12m6ygHHgO8ng9ZYH
H0ahSFWiK5iNmMeTzc30duEMTHHhD27a51jqGIUCeymL9zF1i2slxu69piVW8PAYfJkRXQpDYlFQ
Nki24vw6U2TjTgdDgu8YRH28dV878UcvgsYJ1mb8OYQoLk0gtUedPkSBkinMVjPS8A6STrAXbN9h
DAuYVseRT/qtpemweXytEdNZxIcbZ9pHsI71L6WNWSjYgBUZlEmWA9Eb0Nh1ti6SHZHK/zPLV2em
4MNeXgnsfh1U297QW/kj9feMUot00pUojI8FvYYcfysRZ0TPMYhWtZm0JiSQf8teuEgyyXatCX4C
sSK7k/27GA3FD9LW/kcGocslm9giF+j4HjJfO/PaBPz3nFbsLlusqmrbReWaB0Uff56ZeMT7Bc5f
iVTEa3vYsxqexQo2P1J/4x51U3166BaBh3porzqY5iaHrW0FEqwAswWhXEP/JlGWFJUt4qZPOObD
aeCKJwr4TlxkjpcJXGg4cQrFrItkPHVvlre8xYmpMI1SbXrW8m72Sw6JdyH92t63yLpFEFftMHTG
51oBODpnBEPkrGA4rpjt7daY7r9Z5AT2zSNW6D1/m5eYZ58YFORuYoMkifef4crZeiOg4zMz9Cer
oOhufgA38HKpPuRhcYCv1R2jaI0MozhTnsHk3zmW3T4HsRclEipHBbtLbyIgUdiOP0vNb1/w8QlM
18i/0TZqzLrFCrUOm8GvJVFYtHbNPfRsjTn3jSqdV7v56+7+6456In5+ARFC6G1d2ccM75Foa+Yl
1k8m476WAEmS5jyl6ZTAH708Tbz50I2BLEypYqGTqMGMNLhgfMI94ncmdRKp1A6cLSHZmZvNpvhU
kOAhsZnNDZCjiOW84iFeSwOuHOYSSQKQiM1WAh5ZvWypQUbpMkjX9VXZ3NiRUIWu3H8P7CEhvrKg
zhyKLw0CQe06zZYQZT89WVSDYy7XeZkB/4fXTj6KGw7zYV4fxAlVTcAcWoKmk88jkl5AdYGN6Msb
lXrDjqbgfGpQvc1AbdII4uIICWZiTKaH05Af1uc30rBSk+wUKuIfnCxcqilQwVRRUS7ITfCZjM81
JrCqsBwNItxsb5qN8enAQBRsW6sDoO7igM17dncoUTNBBGq1CN515XaJzx/4I2Fd1HWO4b10frkr
02m85P16XyRTP/D0XnS5g/5J2S6nMhQ8VlnAIcZWH8epSl9DIXlyqoud6jDBJJm+Dug/fdn9eOXR
a0QijSPll5CHA1UVCq542ssGwCa+7zmxMO8rhybYtrt0g0ARbr/grhqM/kDbsxDdA70TeM1Zs3jk
EGfrVA5lD/XCawjv0xtctf8HChHUmgrMAvMbd9gAvgjL1AuOWykPIAVIqWVjm+6IqK075gG6f1bE
lDqmLq0HRm3c2fiAIJiO7Zte66hQMXweJnNqByI3ieutgz4JcifuahyDVmYaxjmo+Eka8yDA9jK1
2d0Q19df6zMcqq+ESwpyQzFQ/I9hZAknlaIQAWxeEROGqEwqLwfhkAJde9eJliZFGsolWQrj3mDj
iaHfJJaJ2ktd4ev10lybdjUwbRekVjZ+rjO08RnZMGyayGpfZ8vMKRLCjhaExVaU5/BMf901U7w6
EiSGy6aJdA3680awEUTPSWNzvND89ONACiyNWqYnlECpjYNJ40kkVsUiil2QgFgrzOLMBopEHuXo
nB6ov39fnGLWVwegbpDtZDGf2LYu10z+EQ42tiiimMZFelTRs99ApCc476yITc+lOiNakn67sMZ1
4wBweJLuL6E8XyrKT5ETzCu9KOykEbHoMykxU3IIYFs/m7NEAXeadnavetbIsdDfrbzvALz0jsjF
jQEWkMIJ0d76BPHm65j3MPAA/T7nxtsgvTf51Z5hjm7mW6I82mKhdvkepltBWVpdgwNA35CTlu6S
j2ya+rz2MJ198p0ogn6pH77eWXYDq6kAfLqh1ZSyORkeOjq9JK1O18qZFSxa0/HZEIemISuhrVZ7
YThatk7UzzHe7MnM9cr5ZHrs572UwpmNHX8uai02oF0K4aqDdxGqDE+bkATfU3Eg4IK0IPPX77rZ
qjEKXXab1T3+QMlrG4s+Tk8+4GwCYqg6NEW7x91jgN4+KvlgMp/6z3g0yF+ea2Kv1CdcwcO0oLSW
tAkrWIGpxcF8bGrUrOXgSHhgwI32zM5YJeaIZHEA8EUIkso9Ig6Vu/xn5VZm3LjvOn3bpOBpOErw
vyG7idJ/GBEaB1muR33/PB7YcyGKModqBslT8tAJS09uG1tqFCK1iDfuJSZjUHUug0BULtoFCwoD
yYtYIMsp8K/1We6ZS36CUNozhO9kobwU85A4hf5duhxkU03H4aehN6aerOvtjLBwgCcouDgK08Uh
cfOUMs5xpjKO+6t9Tx3bcROKHC1pVCePRAZ5yn2JOJyI6GVukG61ueRynY/TzdK1i2rdRSlCrqs3
38iSZUWkQxW3GA7JZl9/o2X3KUJA42pLa9uyfxoyOKNWAn57Knw9T5C1GeHLSjpkDgTZB9mTlMJ+
LacNxbe1J+WFpehJkWwVBqJztMYekNOwAtiDn5W7cJfjc7zp4cu34nH2tErQrmLiEHj0tcXDym15
rSWtMwjjMCmJRZfs25+bDONj2aU2u6fVGTHQ+w58OJH0gFKJtEEQZyoh0tndiZXJVqqJWyC73Yia
SfgFqW2W4g0OdR/RwliwgPFkUUPIOC3vusPrTXMbOHffdFmlzdt6F8zl06plGeDgPsWlSCZjx0hl
A6ueYLINf4VjxFkkBZk1BEdkMfJZIuiI4komV6hFooJqvfqsNeElg/3MEhc8OuIZq9gta5Ts7a9r
T4OQLicy6lDyvtjgxZPgNM0fWbM2mXI8H50RZrhNTrEnHFPgBz+eyx6J0TgtRbCcUidmdO9dhXdz
Y359F/EupHg8xKoWKq8kNBKMx6BpajWWcQmybE7V3Ue+5s65YUjng2+CjEVPbE0VepWEpOFHaa14
pGckaQuLoRHahXr2b79ZKSY3nmlX2UC8dZUxLGYUCOfETaNC927XJkU3cCkoBjR3uhIXfx6ghTFY
z6gEoASgxRhk96v2gFTt7m0ytAHUyIBXeFxLtyMeb/yJ+X2JHfiyT/qALepcILM4SV0a6mmHyWaq
uvII8Km6IM85LaGU0l2kjiZNGBqrvgIJ2Z7HlKQcG34Rg7aG8pm50A/DJYhzAVSBqx90ISf7DzAn
TJJx3D0KIc8rSIMg/FXXGQOezBV9R9mFc7tMZ/QwhVgZnzQjBf4N6ke3stFLyMRUzEJHN5F6iIgt
MgcA6hTxb7uv2wV7duRfq6qZYULa7U+AtvnalTyuQ9UwCg62f0/GT67GSdQ53BbSVoS7HlBNCRCr
5NlINUxoP82wBULpIw==
`protect end_protected
