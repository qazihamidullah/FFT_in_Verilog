-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
VuKDvEsyxWvVEnYAtjzFaPoLFx3Xc/2Pbi5D+KWmWn73CzAf+zAqH3aa6v9BeYKJ022XQV5I6LB0
sQud7y5eEhQuqGEJ0mKClDZBLYdkQ5AfoJKoM5+KBWjw8oNjMghDN6uKR0Q8vkVvoQvc+okNRfMf
XMwpDHjwMFzXdCbqFBYwHZcl9HD0no4kX/sIbMhQOoijkJGaTXduQ3NNaw9q4DwHTAOFXuC2v1uF
a18ZJCi9I6uVBC7uiV7o6ZsuXxz4qukXmkeROI+oFcHSto/QO0NE/uu8BrMozfDT4Q52AHEx+Ui9
lA7wEauE7xXiEaaJ/Ub5g9tKpwlwCLiNClQZkw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28512)
`protect data_block
MoPNx4trlgjGh/owW/thwj3Zp/IgGXHbCBY56pa335S7rCa6TOAWG7VOObdZpzCXtAuQr4GDNDvz
nDyOiM1G5Cy8G1KJ8n5zuh1s2UYMSfNzvFtO4LQe9bBM7GSL8X5AC9CsgJa8RPfJeT2x5tcywJ6/
d677LBrGNBaQB6i4B8nftH9GZftvS9nVX3knp/lBcWx9h9q3BEqkMrtrb9ivN2eF6cpYUHUDWJxn
ZL9Y+NayCQH2W+eUqh+nXDF11ozpjyVhkdQAC9A3862DwkMd3DGxvT34vKSf3S4rTVPfD2YslY1r
2gxWWfEP4clQppyNBhT7x3VXk7jaVlGh4XgqJOGI6kakMBk6ycg5TknJSmV7TBR22ApZYcC8JDt6
Ha2Yrt9rktcRJXLQBoseohHkz9Fmg7Gk7HslRBGOvnPU5oCraimrDUl5VInLy+cDQN6v7YCZWhq/
dn+v5Ja2TZQEt1Teub0lqYx5Q4e/qEskHFcBbXfe8sYiRqSzeoupx6L0l9hlZIC5FAY45YzESI3u
hYTQTSzb8eGBweAG7BmDeEzyBI5mEjFBm3hLUourVNlrnJSupLx1HDVLiztfEXZtuE42+stwwegL
Sj7jcIO9iDqkRXdHdWbZSMEcsh+LYgBl4GnxFKuOMpVaYRqZz+QrnTLdcE9VDe2Ep5kMaKCnRoBX
LOHRPUINDw40qioXmJExuLbn4urjYYVgJIs8ScE2JA+FbofBPu3u0h06anwlKOkyvWxU6tMk6bZI
u+RI8ajAFoYMrZytGJ5BwQkgiAJoVwoJeJQLoiMP8LThncOWPsirmtdIpuGNuvkvzhfhfTCHagJV
COO7jhpx/e311B5478RdPZy62CxEmCiYtt+4T+nmWtBNnKNrTFn6qF5HRRN2c4EHXcBNCJvfN5Ed
ET1LNiwNIdxlCOcTiKguTEoQemC0CNG+IBSGJRN+HNoCEyXjTIz+jXbi4/OEjPWVvtVzI/vZQy8h
1C0cSvtqhWTJHGaGDQ6GjP4doY+eRAH27O62iX+vFuYRE0inECNAnwrx3597d0+QIkfVAGOmibJ8
rFAtZMlXP2lYpP0hCDp9IhZv8B1yfIVEyvVofg34yI+YKQPEsX/yR3axWUEZQqQTkvxXrVrWRdaB
4qlwd2bMSHgaXWX6AMd2zUFfhkmiRUpmzRT5CWMLXzgMQGAcJm051UVuyTXx/mJlCF5d5mNCHmTF
oGlbvqGo/XxG32UNq2hDrd+ZujwyzH+tnfxkDG2PIF48TJxJnyvhQt8ZYfnmg5mEXxhz5QPqhCvc
56kBRKd+tg+PBYVcMrsPQVuXAGZx7c8KHq56zHP5+3E7PK/0IYNq7BiztlW4yqbGi7VwkqyMcmxP
H+V49tS/L/JgPV5yHTGSfohdxDuWaHmJt5LmIAHlimxka1lV3BJ7t5JVK1ZuTVhB+/HsPt7Ii+7P
SqTdigcQRI5eow+0w+lonCvmO+eQ7qjCjf484Zp0I9yR4XPQVLOQSj/IlavJOAm8dwSJgdwgFTnO
lVDmiQamNw/Jsw8GEGee+W90lh+PbjGWqlNeVnh8UZFju6uHogmQs599NRg7AjLrSsSkOeeP3v80
w5Gy6DmvTLr9zQ9PBHt5GL/vutUQS3ExrfkaTaDYTagxLJ6zeR+WykanzVxxpzXz9Un+t1uplcdQ
Eo37rUyHgsMCnX1UOM05eN1hVfSSGYNmM0ZWM6NlVCoC2IRVlIrXPDMTuOHSnudg0LpBJTm3EgmK
YtWoNWZgK4FTKI9eONwhUKbs59ucjZ6kywg/+4SFGCS6FNsdp9re5TBjVFOBn7ZQx0OxVzRqz43d
Om6UGrDt4kdkm4WaDQNgty2nvcvAz8TDJk+B7wDLdjdl1HZSlTF5k/XJqfhd7GxUvqWhLzOAhTxZ
NDUaPE3qC56yaF1XQQDofaInNCELYraf+GhgPFiTbeaNCbSF4vreA/iZfvJcaOIg1O1J7xQ9EJVs
0Qwwdrrm8azXuj/9QbD2AYorNwz1Ee0zDctFjMhL3ZvzeodTgXIbiGTl6D5m4OtJPIufRkA8lN++
V59vqn/7G4VM8zZHhNFVYr2lrQVzyiBwiExqHT/2o9wmIhxmDOFnxkchIqF/mm1zQtpiYQdrMtMn
pfjEQnU0dTkknoDDn4Nse66VA7c9yrlCHNcoOnxyk32vyBcmAPfMIL6YIqjgbOVLSjs6fB+Nn1Yd
VjjH0XurBLfipSyu+Jl3e+mU46w9pz7hWvCVLBODekc2Auzblfxocx4NWvFOiZK8vhOndeIaAHyu
iFPEOKUy/bXbJRRQEaOaMGlYqEqipT+k3ewnsplE/zm5aNvKzDrjA/bFA//L1uNW7vPlSGUS6eNC
WZHwiQYZuDkhE47VgTu7B+/hsf+z1K7S662PGo9Lumlsq3C+QE67xZN3vK445pVyBcu8BQYSoFdP
BTi+SHGFq+mlKLUEe4bkKrOrdVGMpLoCgdhcwne9MekoTleghKN5bvx0/q0uLhWGs/yFeKU9f354
QFUNcCT/iwgaKMxj8Ai/aLOt5s9AdMS0HyV+UdABX/7aDXEBApr0CM5Mx6QeuxPgouroS/wYdld7
y2Vk23ZvM3Xrdo9vre6b6+u/4OT9AobbbY/U36/59rfKH902NTWmseMpaIfgdd5/ZooQ+pcy52tC
kdfNIOMOpbBwMpFD5WyB78I3nIXKlktitudYx6U5Z2/r8e6W5KywZSo7eGcn+Hgwdw8K6wt3doeA
aQ1qBLCBjZ9Y38TUh7IA2yyVKlydRzGOdu1shlGqeGxl0h1LCAkKf87BKXy6y3xAwtCwxx2o3cBy
HTNUwzAxzkrbsSAacdAlOE5fHTkjNO/5MH59MphYNoDPSjoQuakxI9QoBMROrwbaMtudtr6f5TrK
gegO/0cQuR1xwCKWDJkuzmA1yZqqbVbUsDB0vrGY3Xn6TC1PrxWVlzS9bw5QtudXaRMUpTL9lvKe
xInV8zB2AzkJvpNNxqUMP4sg+MI7c5XuaA7MWgs8uHgkfuMgHRNrmBFgkjShAroX3SPVCOd7GYau
bxcSn4B38PVfnjpDmZZT0oyf/Cea3XxasOTb2T1HBS7dlGFBnv6N+2pJ2GTWrdAdnR/Mr8YApJUE
36Vcm2pTzVpoHflNwrNM3UhDmcFay/bGyd7QJNGHz8qCCwjme5LSYzoexEopNuUOFveQKD6C5u7c
Q92LDInjBgr+cddI1EPXrUcrceHtimeuwi+/DWhlmUmsu1jIQJ2TXsV1ky/mJPJGy/6b1ZzZgIds
8ZXG9xj8S3vcwBS86ftjokMHRKDUDobeQEtqna2n8rRe1SfdhX4YSuYfYdCxRwwaw81CYJ2MAExt
JiDIaMk46I+XTzmTNO+M/Z0LNz69iNH/HFYtoC90J8NehPxlZ44l06fS6+R1a8VzSBrL0oN8hETa
BLtQ6uekY9jczeaCSNiOyo7WMb5PwiGPRu2zMwZna/mOnzjcLI4XyRDu9yw9KamLHhSyw8QmbSYg
ZqYyTujnUaB7TvdHcghenCPbenT5GNeuv5Z+8mfLQmRruuZ21zSZY+Qnn9ouN1DR14jthxCJ8T6e
cTLxACFerB+pg4fZUDkxnxuBsNHdwCqpbX8CfYyfQ8ieKmdUBRH+0LWhd1J3au5AUrvEwDNxN8n9
apS3yrXWeSayKdcdgwJGyDU6pE1wMbh+AaYoSTX1IQfbc8Zti1u013wR2K9TNBm6CBg9lBJq8UN4
OBBe1odMNXn+N5yTW76EAegqRiMUc4zYTZ9IABA43QwDyk+yFuCIaYBEuTR8+anQ6QhwpHOtUE7F
EoOTR4h6sFlLo+mG6vThsqS/uJEt4TnocyopGIaT8iQX/ajocQCuXhWkYBwirIAWF8Mpy/x7oxzw
SrUlkWCY3xn7Z9lnztGK8QvZuvYuvCXDlGcWocEhuA+rwD26UYcExLHrO9ZFSNJqwAdX+XItCCld
QE/bL6Xc1dtGlfKSP69Alp4GrcRcQiS28T0g2pIdn4Ap8C5rrIAtr7uIrKVKyEjNnnxiuVtTT/qj
aSEGjNsJ8RRzQCRwH8xhF61BHtDfveKH/bnl3+UU58X8A6BcmT7SYKdtModBzBCkl8tzyAolhfPH
UW4adYbGL14cfXcouu5mAvADHBzVn+tMGy+WN8jT1I0W8VxKoBovEZjirrNoTtvyyHrodSbglXsz
rCZeW8KOoLt5KR1wcK8GJ49TFc/V7HZSJmy0D6pMmhj9Pdhrz0hW/WP49E+UBOUB3kE4Av4N7GCS
NM5l0HtywNvCZbYSlbgbPjWGwoQAXs+LX8EVsGETuvH1NE3xAJRy4+Gno+Nz+7Pem7xig1r4Gk/Z
4OpxViBwyEHcQEdnEXTqtGfFf9/0vDfkotS/SVMWtk841u9tQYP+LdXXo/vf9/q9SxjNSDFUPQ0A
Aci9QX/OWRh34WO3l2XlXVkr0rj174mdh4hGKAk9FS9pl06hXaYVHniHjNh/erEA3JxN5mlYRKH2
plI3nkxndT5dbNJj9l6WmDYXgfKvbEuSuYcnorP2xDs8IpjLs4ybh8FJJeXHo56Tv51od9MLRGvK
JsLOjbvm6u4CX3zJRn8e4bOPPNxmqG1QfpZggDNot0aWr4HdnGMaOAQ5HTWBS/oN5JEoLe+CjO7Q
YMMTtz9QYIzrkQPjOMp8a7dcMncdwjPsiOoz7NyJwlUJZmNHwdPkd9uANLQyuaygPbW6JUNykdvl
xN82685UcnCdJ4Vvkx2xt3gfSm7rbiWbkoJjDxoM7OrKs4DoCdFXDqNyQTQXt8+0gXNt+p3nKNdP
T87qv3mSMkkw4HVG33cFG9iWAE7D9+snqThE7rqs91BpGmYVHGeSgwcntEI96YbhdshmWnwoD6wn
1OqBQc2zAVWqu+kYfSMksv34VKoD72PEjCKAB7EA3NLMOuxwFcT1iiEXpY3bUm9UE3xIEYxIxJV0
hTfvL6T1pbfPdim1W3jUv7GpCCE04W0ti2WGZVeALOrWfBk3mcQNQq/PgD+4eK62NkEc0udKt8Mz
MmKlgIiq2wlOkZH+o6xgV0S4DKwIF7dEMC8mZGQvliUlm1j5ZMrLlrhvlYpurZ6tBZlgJ9392y/Q
BlZDBrjBt04prMjTliijMywMsOBD4MJkZSo7CVAcJKbzGTvbpoz/5wBKbRd4M7eG8PsH0EfE0CY/
ge9NwqW906zgGaDrWAMbJRHKFGr2BC8QH0kdNTSvSwBY3c6T38FwI51hYLr5hcAugOdZuMxtpFXb
l7d1BC9Kg/4JDYsuHyY234SUSsgEbUWQcdQX//l0JS82Hjkq77CWrmRRoe/1Z/FwlEZ/1991VRwL
H2C65J0cYXCfgdN9u/EiWqnRj9ubJe3TEpZ6wZhRts/08iwPOE1d6G8+M/y9GLXVyEbHlvuQCacN
xzbv3BmMx+mVRRSBXFnvdhEEPFW00h20pVKR2qwOjeyKZBhMSRDlcNhGi3YkM7/67rDQ4oVvSijJ
TZ/IyEHOCwtaSKw4rswaTR/SC9Cu1POj77Coy7+rI/fMTG1h97iS5xVJLRN+J26Ix1wgiDc3sN/G
9nithee5AsIM3BoePj2DyeKQGtpM/cXWKc34OE0OWyIVRgU2CwDuOcMdbJnE17LNhClGonqkWIdN
qE0E3+ciyXYGg2rb04QaKm4zlsU1ZC5LLc6u5pHsuuFn9AyqfCF7p21xn8oT3xn0BWvy17q+HMCA
T89SnNaWGVhitg5iAJ5jfrmmS0VyPGeHUatUWIC7GaaWZPklCQUWvMAjnSZL1QCzip/14NAaF9d7
IC9XyI+9+Yhv1aQr1G8qaShIbNAEGak82MA5FcCMZhdr2RVdqLcP2ZGH+CLGQuvSXpUl+qU7vlt7
ujTZZIklxn2hG3D4FQs60zQoYpxjlxRw2hpb1UP2vEuyISiNvC/ud+fIhXW6UXGt/P5DBcwjAzfz
3U+bO4ccoTbmVB7mKurax0AYgYNpKzkzTQBvnJwNZR7A68SRweJWP4eSOS1UDCga8JgpUyAoo4c2
9azi9A0CN7Ya9VBTI1VpIC0/r8F96tsmZKo3PeGUBw/wqrP7IEWrBacILPByX3SQGraYd1uba4EI
+7a+GPg2tyP+kr44VdloiYAHpMU5qB63p+UnKEgO9pivkxIVeWWBg+XmrjKBFfJpKf0vIjx52qrT
tGTW1nxBHPlSBhNyMm0Kwjc0pC6tRtAcp8CFnSxbOaWpcKsfqXL343/0lKTdNu4AHmf5orFDNNj2
yV7iUI7ELpHdp0qB9zK8cvpwAN434w+FPBI9QiD6V0kkYZ1CaHYutO2jsxTNSFk0R5rryWHrSBXi
3QGGDT5FY36OkJfZ0Fv3oYXaQVxaLSeGDMCpn7pzUqZqH+PfP7hfEZgx7BXhKpORoLkB7J8s8g9X
XI5ihIOtmO+mpVnm923e9HJ5zdwjxGTxAdrqg7VZJqUnutcgG8R3d4eAqnIpEuhVHfLMuIuTgXkB
A24WkmpBkEb41b33VCU9LGf7qBSzFVynuGB6Q0F/LUVNgoFKjoGhTmggnyucMM52wxSd4PlUYK1N
CppmJpG6cge6x0sKXj8aWbL7a6dcizrr9ioaI16MrlGLWAa/zwPoLbNqliQn+GeUA53G/aDA7VRC
7QITFVhOEtePqvXJyAGnR1fO2EFWf19lQ0vfzPUFRqugf/Y6G56vuyHzDyc2XgMWBIdX5CfNHWPV
uyqWYqLXmRFbSiSFQjGoB9pacTB7fT625CuFqiqL8AqNng9zStGRNE6aupmSB9uXvj7CmpYymgVq
Ax7LtVGBPeNeMYpfxUSMsxq7ol/drdMiRcR/RRLnID8zjPnrysTlufJOgRl5esKXG8Ieb65uOazS
mP5hEnMniAK3B5N0LWOux1+ezZgTfxDhBi+0Eyx3t8r7I0F0Wz6LJVX3m0CUYsAWoMBMCWAhrRPp
laPr26a+Gg7EiDVnxxiaC8aZEeaStKCXTFQmnI6NWz8HtZkCXvuoc6hZ7+TRcFKJOK8u1WqgQ+xt
m5NQgA6a5LkPMvEeuIgKl7er1D2cEjbkoHFPFB4JBE8QdkB7EaBbfYZJl/GGiDfn3vfXVGkTPP63
uwgLW1gHBBu2JYo69Mjy1NEfpl7/7B/idh+WcwpRXkoZP3V6t/RfwBiCMMCOkakRfoVSl9ZttwbR
30/XWiD8LZ0658QNlzliwJZ/JtNd+CT6ZLCLH2UsI8QmWXwILqyIl5ZhHZT9ZwzVpyGNpf3oeTIb
Kvqtj/U4qnGxI85agKsEAlcJId0aRvdo44dtiXaDbMHhQDIYzWWoqj7Qud3pY46ba3fNVb3m/Icv
W+I8hCej0n+z40EXbEEtYsrwFCBAKla9pGslAmCjIEQL8DZ9mAyEsHRszxGFXMxSh2ezvEWBDmu2
r6qVvWV9PfeRSwcFh6vza6Je4NsiEKeuLN1YryPvKNEZDULvTRMBzipGtDXBUoos/FFptu9nzLp5
OFei5ewKvzOr4Kdd72fJJiMElE95o9yhtfSaFNkUeZ4JCgZIQon3LmQkFBnEemjp8NbX92kmYyQg
WK7ysYMmkbo40qD4FnXiAzAaM+M4BTXTtSXzy3lcqcS8bHtxMyNGpdufORFqnpfueaK1zGmhrJR5
+4XAyUyanen421sF1CQ/d9lWNwi190nlTuLuN56UcyGf30NqW4Jz25H5IJHXsqnOItTebSm0zdM3
OAD58dE62hxnrqLFzKsgUFjlDrpQ+5xSNVnhkMawX0V7L+YLmfMYDkJTCIms2BEjbUqKZ3pYpDYG
xijGgtgTajWUAtNZwIL3W6n+Zyg4qOfpq6ZJMSpgLT/L2VxDaxX3ijv4X4UXM5gItKMC2zqlircS
lhCAxXpm9OuydiAfRGyccbo9B1i7Na4Dva3qVyhHNsJ5ijgIVrHFYXkjFG8NWJ21Xrmh3icXop1O
6VxoRhD2pz9lvmWLuNWPwRjYUUJXa9u6mN1TG2oAPFgUnVh7RGndPQuzK12/prNyGzsSQJK5q8jX
QnjTmcNOtj4G7ImpI8JJNOQ+T4p9IdU/0JTs1r/PNpr9DyvXSD/7Ud2XJvD6XMuDQwfmHgj4PaKh
ecLItI2F9OgxDG/KeVgR5Izq5P7aHMEMO/bz+ZvKFmJ8FnipyHJ6fhnoVxM6C4l7I4S73fNXG8xg
CgTs1Qrui7cagXhGQNdW9cJZA97xKvGQzETIeMEGoGgsN+ACxqdN8zsb7Deh30gt4WoIgQdy+OB4
vN/DWxtJIigVXfpIOz+r/46fzWWCaEE5UAElFVI64T5DD59oe2htvlzLpbafOo+TqtYQahx0i37d
NVnPiIRBYW11fhtM+tS7P0AT161HNcj8hT8mbWLGxK7oOceB+DJlquUGTtqcjyvP2Mg8kRMiV+Lx
VGx4c1Lyvk9g8IrIGD16dheOeRa1qLQnw8HZ9mLqQNqO9dQMFGMivWEIIa3Rbl/5OTx6y09vaOQs
i47kB1e3+SdgHw5WTchVmhG+Y7w1b2xlf6J6BtoRHsV32g82+Dr29yHZf5lSQGjYqe8Kt9GGdNOK
qhHtsyT5b4emszRkHMO1+GHQLIH38Dx6N8Wty5aKbjbL+ccdCzYH2aif7ywomJGJQY71jvu2FQJG
YRDNrfURcQmwVqHYikjNWSBcH30YUV3W8dgITDcudWV9H9vSMbVcn3uH5w60IhUyRwE1mhzk8KdF
i2WWczuehYTa9qAwtzDe7BpxegijUjjiB4rGBY3Bdm4gX2v5KO8Rh/mkpGiEha4+4Hg+wHGLzlM/
QP0xQnqa63Qu38vu8D7mtIUDuJs7EmENGiAl4bh3FtPG+1wNtNcNx8P3xAYAyVMwOu0mgE4/gz1P
booxm/edLQTq1q6180EjLZbdv31W63g1SCNY0Sc/VScULJ4qXOPOnL9eBSkkNEOPaRAZTxbU9WWe
b9NE3DgL8+oVK7xOdDl6zVb+MGuNmvSz2oWpMkkjbzNxTUBofTmio4uQR7mMqgEq4LeWkpm3zgrr
rzTQkRTm3ui212i3LYvkjgIQpbrTY8DUsUdCv7KSJE3iQ01r6P7RgZdGNJXGOkXW+sgJVuwvNEdl
Pn+gkZAvbxeRS2CZa70YoymGAQ21ugKUAY3M9hGGL7l/Atot7SeZETZZiR4mbbpf7ClkjSL3kFWY
JdlqBjeVHxzLSziVlpRvI1sZ3aZ2Y+HS6ugNTaT090j+j9pgvos/CsW7YIomg2MNy7xGOeCsoS6R
RkAvovg2dxoWVSSd40gM9bCEE8nKBuhin4gWPOQzPydn3rvs/Nrg2CSFr9CYAONO6LQpivLNW1Lw
PmkdVgaeHOvrJym8eQ/PU8FTBd8TSCQ5qCYBNXf7bQ8iKxfKXa26k5sE3NhazOdhen81aN2t94rN
O8mds/f9Z6zTrXAPunREqqLC02KMwFhYkEkj/qjmJyHfsY731HGxHRB/FO/PIMufoFuGDuarQJCJ
YM9Nm7iiq6iM0hyRWR8UFSR+HplcY91coT2Gn/NEgoKu4uPWy2OkuOAuiHwQ5lVYYl8Vk4SAx1e0
9zGTBqssfZ8WJYkT2aeyv5ndfvTlsBZjlu2E2dgvmpyjVXBCB8E6icuB/A8PmrPihqjJzYEL2wLs
jzDgonVf0iS1bM8Gxb1I8mnm6doOUPwuqxdAVQaXrE7jneBWn5Fnc0BXLdAea8tSpkwYk1SWGBPb
pfcworTR1DPw6nTVr5ijFlegVImqbj8VTH+/QUlVcyR5B5Sl2s/uam1IjLi4F7hzTvoIs8vH6IZh
6FZit4miHzwkC7XDa+XddNzs/rk8bacPGG7HvU5VqxOVTnYe0t1+9OWlaomnjsAsCG9uRqAQuWza
F2NbNx4uLpH+bTTuAas5tLc7aeWNzyo/IQyuXB+LmYAyYKgj32VDhWyMBBvLkc4+/XdWAxVSivCm
VT67WjGBBcI3tmWmTur+aoLK3kf7arNVKcYTKglaww+BTCYiCWYiUEHPed5GSt7jcWITCbxGTdxC
YDRuXuFKlO8YXd6mX1lR4Aw9xtVnG1zkdrCO0WGascfrww+oH3mpHR5EPlcaoudmJ2cPdgIjmL5b
qduXsI3GC5OXS28fyuoox0qKS7LxFSevCKAKWLYizYNoq3IGUkpd1S6MOffDwHMjyVfIgjJWfcIt
Wezi1JKgpnpXAAa0n71tKCCBY/IbxGBzGd0O/3kLGIzK7T+SrZfG4169I+ocw1XZRlNyLfbbXwYA
A5V5D7JaRlF8cWYqjNwCyZoaZcUtohOdOh3/G61d4aiU6Kwm8cvxYKniOUfm1yCA4ocp15lW120d
mMaEqbk42oImKpkXYWuzqGH90yRoqMIiGWWF12i/PXkeUnEI5pz9a0fg19xt3dmhOIkSdvxITZtI
zDWFBnlEKLP2rMjin4k4vMEnxz9xtNeqYftFNQm9Zl8aO7G5qqS4sPGQavgrLsEWWx8rhF70oNBa
ygvruDIfOVw9IqFhR7I6a/7p+fkovKQg6Pjql8DisI7xK9tgVN6/wZKUonJ04exXA1qryXSuKAH1
aTKw+7Sb73iXL4YXD7Pzd3S20morfI7fwGOBFQFgSPejfuJl2/KeDYmTdpnq5J4YMbuYecYOTr+v
+lpzPJFpy6DHPqrHvECYvX0cE51nwwEg2xWS89ZmbQSdcR/NCneioCVISRI6xVnx2Q5lWbW857FG
b2gJF9Ol1MgBPyRSlPvQaxP4UlfxyWIWAadpkXr5xpPZpGozW8UCaE9gXchPk5pp3kLGYs8j9VM4
rTQOrX38FyNSmPRK+T2WgeA5NPnMK66NzA/4NKZkGvD9Pa9IEuqCrHarH6htXGnqhBxD6GuXHDoS
Z4n+XALC5zwVV2PTWDOo9oQ2GV0T7IkL2HcPki2KYchv59INpHtM3jnt6Mt4UpxXOF6gAD+JFNJN
1KpCB/hn/aaj53P+/nmfCMMlEleND8cwP9zUHGOsGy8zlqzJQwjxB2XrSAoGk1QdpTjXmLHxAxi3
Wjud67devuISfU5wIS7ml4Avn3pCbQo7GSMg/SWadb1f4IxfZMUU6WZfZsBpG4rZJTmEV4Qr3H8W
fR99CGK4Wf4DFfCckRvM/5hxjNtbuA1wo27HWOnrHjWY1HeQlwcwoFiKv/l5ca7OrCJJ2WAwGQIy
knfvzF+eOzaemF+oU8Q3g7S8M93XLfK9ZTQwGXuZxs7DmSc/YoPnd+bt2/QT5ElnJClFBpaYBW0c
9nb1Xgd7avjTvD+4+dRqTuusmz/eGozWpXh/tHitVXcyXsoDM2/8q1BwP4B17gkwBDWO7XKYhhf/
2D3+ahYkcQFWg0EYYDlp9AkfD/doDCEZbxmFHioUPiUyGYFg0mnQRlwe91UAFj1RTCH761ykwtA2
VfA53Ah75UAqJEs+f8XeuCd4AgH7bkh/xDIfxXd3bNSiP4pQfZjzDuIhQeTmkaNymnlaPuGVINai
mvhvFEmMnTOaJv18R0Cz2koHhL+m8D03Q5OFwXsJxpbNylVco1hqCnhxCuc+ox53BdDu6NuRH/V1
URm+jI2474de3vaKoVxEAWWOje3zVqXgrH62j1SaEelFavYuWxaTS6ayLqBc6z+FL0W4+9p0hJ5w
LUvIj+mfWrwTqy1bJJ67XpdiZPSDo2AQscRuJIdfPEYTWd7XcLBKaqYxsNr069GjdupdpX+1GW+z
ZHWtSRIbaKAdJGfQgeP+B8Q6ZN9XaWhhHSNrrJjoPkJtN5/Dzl2ebAMLSL+VTB/6wFD3u4+By+Bu
SqhVtUQ7hvqJbPXsz5sEVGekRyExUYtLZYfuS565DdyrAb5GQ6jv3RPVRRvpV0ks9zBNwXf6fNue
d4J4mw71OeU2FCMknsyZnUOQjVDhRDoqz5qdvl6soXGI3RtqjLC8q/K20qkUMRFGjd71js2uZaEI
Cz92DCjDHpPTKWVMsWvTjBtts3jqhFw+HE1WRg9kZ1VswxIpgLyOxesAmrCZofFAjBVfTR5WQwBp
DjYCUJt5nDSstLSOWUpKQW3kuWEDwtDfBvaZ6SgSILCz6yo6mhs6IaH+eF3F70pwOffoYVf/iqqe
g5MdorlhDatRsp0gfcVIasIJNeOxHcVKmrGTS7OBWGBH/hIkOPbD3BqxS4e7C1nnIaFxJXSYLUqQ
ps7jt+SOajm8ghWWvPxkbmkiPszAPRcHvmN0bxLjNapztUxE5HXtV5C0YcW0WWyNJupPY9m9Uv9A
cz4BLvh0v31dMkKDbYAQKV+CYNDxAz/Jxqz+6+IljHQjfAweytiVfgUzKfnJdFu8mYx7jJHd2kVH
CTquEzaWJTJGs4FOnupwIcblNXAztq3p4eqfAM6/F3xpjckrkKFvrgup7Cx++DqsW5O/Rn/Ah0pQ
0FyBmntFmREQMjxYycNq/bGECZrgF8ZNjNnT9vgRMQhknC1XkvF5Sw6A6Wc7odyOstAc5o2CmTyD
tf5PkGLczdlBOdD1M5O11mFppuO4EKYMGv8ol8eHbDkCtcVV6KbYfkuZq1+XsRFte5AIQxxJqR2X
y2WqW/IGdxHBde6v5sHwcKErQLR6FP27Bu1f2y7rJ5PrvdkKk2SFwXtOWUsGA8nQcxFyj54XglLV
at7io+Q2ccQq0fb0jnNk7NaAYDo7qq6YrC3tdkkaAvwqmCkD7ETPE23dTaBQn1kWfCS+Sx3LRRvu
SJWpY1/e/TpPQX9oem1ROQavH78EuvmO5X4Cwmvbr3CVyW2Jy8CiuogMXYzg1bdRX0EULpxeDPuj
AuE5MGsZWpXvB5vDHbRan30UwmVGy+67Cy1f2GOhGepUhefROmnvIIOWmWbTqAwjfPn8CHyYlyog
Hzu5PWiv4trRqFVqJwVpmjMXzC72c+gd9UeTijH7vwcmWe0l4IhHtjZXlblut4RDs3yDxswqqvIV
psK4nb2saFK/2GJHFTSXV+QqxfZ1oazwlMbAA2jhGHbSXsbaJzabqRkAMXTq7K4GRd4dozH1BsU8
Yq+qEbYZ4QT20w0loMsuGSLyVvQaVBFcbNT8emPRRDpU2RMb2x7MhZFP7EPbAJtE6hhfSe4g8IaS
BZgCuJjqHcQeUKPWjq0na0Qz+IGRjZ4mxiewohHVu/yS89JUnMPeuMdXUgAxxDp3HpkVwYTcMBXp
PDDq/e83M5oh5Jgx5oGc6m1mmB1WGtEz/0BegFTKOHRxVPmlFZavB9vzgaz6khnZ95T0R8oNG6mZ
4nWSWbXv5RgNHUJvNMf0BoGtCxVNgUwVtWOAtYegBL27rKINjfq94WcbAH/YD62AvbB6WCosSGxe
slvkM7arnubQYOZMuFdnN8DbH8jVYjk8ZAyRDRp3NLHR6jce+kfjGdyYGrOH8DB8fwoU2tUrQziU
e+thWhAi488dAXlJ6K7XBI6dxYONA8ZEerpaf9NtIOHmX4H5J/k40ZeKtY9eUL+aT961z/4I8n5j
MyyudFNiFdD2qdlFSdMZDzR54VqVeBrN90friYZC8zeH8KC9TDNy5NVE1glIm/WErxm8HdiA0Ixp
FDepFpyrTD0Yb2RJhFBfYrQo1jI2bv+HrirUfy9DEEWaov3Mg4pea1Gse4zxeGGcMyY9JSSDZqIi
J7YLVfUkc5vVB6gwPhU/InOabI/HNtQjqmeJz4y426W9LbvpsXltWBYi8bovIypOvoAzxxI2De1a
AQ1S7TTiyCLwsRj6BzrJPOXG4Eh4ttHr9mEtiP45QEAiIxkb0HWn5kmUau+rlVqECnRLBSz1aRKk
fTFrTZw7kLWUTnK0ifISDS6soUR692G28e4/u5d6QZxYSNO/im+siKghqck7tN2et6MbguTgMejk
5S95jagkP+23eFHETYiL9M97PUiV4KGsD77ycvdnTjB7fuK3g/qYpddv84vHxFnTjn76gGowAviJ
+QWkIjb78k6k9EGARck2+lyxRfgJHU3IiguO/XnxXzrxX2UAaJbBSBfuuXF0DS7Bjrfvd4+EuO0j
27wnCzN2v9JJvKpCXv3vJvWgmP3Wy8jAgjwlzzxFZWJ0L+YnwHl9g8l4LIf77gQ5B07nauKVot8P
nrapa2/InuELrI+OJvXgIIM9BvPjXljk+6h1aP9EcY1p/Ft+QlvNtSU63TjbQ5Dkai8qAlsXC/U5
1khf+8Bhd9hsrAdTi/6QOKllxMnnLJBXQSugKUsWUQ6blM2djajJuQ2SiFvYc4E/mpDrMG6zuZKv
QBC68IeUmKLrWjQ72ey4ZC2EQju22xzIOSJG6reT8joVLRjZm5DuXvcAXbWZt0qN3D5iagqVU1ql
iG9b/+K2wIvaMiqYEYgmKuntjszsKqHfWZosPraABgYNtKPwoTCkBQ62EPS7g57ZktciOFK92QGK
V30+m3nRn7T6GbrXZTqQnvcI9aQEoN9WZm7HsLJxP2Zbx3qte6DGTusXwp0+LOgG18+BM7VmYLaA
nuOh7xiBvc5cggJLC5IRHJRn1Tm3V73P26rvj0O6cgurmGVkHmw1GgQ3wrd7whUndwQYajSH0ZpB
EZDCa+xxrgLhiSpE0tvqvCBAPoUDkJbRRDELAvRK5cld3IC4CK2gmZeY95UD7/lYYJXCkyfHQAA8
R8UbIdDdq1plCU/j8NwG8GHg8TypaseG0ipvujpSmaa/PyJ23SuBPxTUr6Q7y/bIoOifXusoGgDn
qEFhVAPih8Yb+2JpiisLLOJ/xkXP64lmm0O+4vfbTn3CLy0l55itCmsrPVT6l82V5t4u+Elxcpi4
QwHtovgktP/QO4w6k24vSW0zCwYA9pnu0+aeACr1rixdMchm6cnCIUbE+Qw0bIQ9Pk3OZiILnFuO
gvtdQLJSFJgLuThxWjI/akDY+DFZie2kHKvd3fewthwo6huSwtngNZqxM/TvYisuQatZ1JsXrJnl
fXkR9e2HcC1pHOx9BMtLHogIDTFztGM1VhUaeOnO9wqsqDFL2e+2s4TAPVrYbp5yjo3JljYxtcd+
p4JMRqfvsJ5Tkxj1upPvunXvVVWAXh0pbbCQXS+nuLHoi+qGaWlCOa+7hPcFPhM1Yg00OinmIoDv
H59JFdLVx8CMQx/uOrWTWz9JGUVsSrnNk6MITjEYNnVlo3M3Q60xTXCgBckc2hWKFSsS2rYXNK85
V40y9qmcVaciOwtwizEZFIhDwmXP4GysK087aLRfxZr5onRG2pq6vgc2WZt1Eh8QvU5EASAFyCxj
PoxujZf736t80O3BQQLnYrRYFo97Iv+1kQ2rdv5MUNPXHC3U/8q0E6TIrI1OejvxsZtRuZg4CxD6
IIp7qcrZdihnB5r/EN7Id/E0A1fow0OJ5+q94oD6CGH6JkQRRiVhoN1C6b79gjJtIRK5diggDxjR
wjsxMlccCtekvh6optRivcJmKEj+ADY97TGjvW1NI43lm3InHCGEkFRxSmz7MVTcqXWpACaxCeEl
dFFTaAq1lvpOSNb0FyQFMSZS0X/ruimT3McDho0BL4RB33K39HSDO6jyCAnU6Ry7HjEH8C3oukcI
yhJVjV0/1uuOiAun2wHnb6h9V7ktEGXousFDJr9xErmcMrHeQ3r7AaV/GtTL6Fom7dKjLHJDY90l
l4Q63C4iIKxty6l0t3sg/AhSgDAcVl6JK9OvDkhE5RazzFvrMdGz8YE/AVQNyx4lTNht5l9no7rf
Z2jEgy57P9jLrubZldhUDlAYVysLlLl2C4xug9SsjSuQJ2z4tEZzKcfERWcr10/lORXw27GZaaO7
Fhf29uqSxcX1PvsxlFD83BE90Y6FTviRKeHekgtJlk3PHvC1sSTSNgexB2eFPCgqR+TEN5OSWZ9Y
V/kEOpxfuP67cLNRDQuc+5rt6qnnBd1siU0wXqYgK0kW8xF/GezcLg70NvZLx4RxIRL4RFtMEPje
ThG+stW+ufgK7c49eQVHdLrXszalQg4ofC4O367gqU63/Uir4YKL+Dg7Nv0n1cRn8l8AwuxFGQfL
OMa18ZsjJtKe7umRrO+2lSWjjdKQXfkhsbIoGbB5731w7c/Xt4rW4NMUlfyFAUxIkgmCg+NGWWna
yx1oki22GoLukMQFJkRHkBBKk47AWk0PdYGNJfw6dLnHeHCHj/+r54XcNNa7/kPUo6MBWOZ9KP5d
XG6EEUo/VyX3dExeUc0Wbc+bUgeF+S8QTfEs3Ur0x5YUmOhWsGRmY81DrAE9y1YObXm/l7Q+w4qc
PPik20Av/SB0GdmeTIcq5N2kQgabVTAaAhEMU4MFV5cwCTNwv6V0icnHYPkCodQI9+YRX+O4kikH
KJlDzdlVK3aaw0GY1At72FUHaBNWIlXLG3L1WEEVUiwEcHqQM3zZfgQkpQ/TA54EZkqDoEzjnE7L
LVWfUv3vrkCuPhsnQtTx9pG/9RyQqGfZPkA9lSqWhHlhq7XU7wQ4+gWSkeE5rwSeEakbA/wP5wOv
idiB0Q/2qLOrymmyYzRtJTo8CN7xdKCTC8c236JwdvhHbqeQ3VHNwb9r5QJRnGYZk3gDMazqib+H
XEzBKU7OHu3m2fVPkGQ1gLHyacrJ14J9E6vChyHDUU1NjLEvkbSARrACOqsf20bxfmhAkExRkDX3
OykR/nJby1+LR2Q5nSH6HDXKv60XWPTD2bYHgUaaXgbCzsM3j4SWs5BP1p/obBY/LZBrM6pMAYjM
FfObKxME06OyF5KrgEhcZvcjUFwkvNyRx7VgGViwPWc/6m9vQMPb92O295muE0yxvxHZEdHfb6mx
lXcr/6cbkfqD4HyFLCAmr30WrlGXwhCUix8JnWTJ45unr1/KLu1ddCj8TqxSYKvXXDHIERX1oEuZ
u4dumf/fWOf+7PwzmXl4ofiVBfeFp5dg9yJxmnXMaEZX7wRnrZChqepYyzYNLRDsF3t1NJUnYuW6
srT7N+U8/xePjF1Rwtljkpoiz4FGp388AfIcoNQND/iUrn9i1nch40iwrzlQ+oDSsaul9rRt1gDo
rh4j0pK+hEciy5/hzaeE9pzFqtS3+2RWyTPHt84WEh6qjy/FX7UKA4fzcHKoM+c4rTKh6VgkQuUm
+KrRWmS69M3V6MlMsYHTDSQqH6qHZB6mbSQnsqpF4OAjfjZCEzRVQNWjZ2J7kkI+a9oeR5DsJHT8
nYvI0z3xxfTosK0yHzC5KJCFY5ENrQmTr0SRSx5dQybeh40yGcX35npUwYvhXescX1ea8KFcBs3i
dtfvVoOiW8wrKXXUgRho7hCtbJBGr6PskzMIzYtw9UetNmDh/Tf7LkNEoOzv6XDUnnrnErDo5I7M
oybmyG7ulkeWfqwPP2mWmtltk435uail7H7KsaA8laUWnFHmrSVkJyRR+OBHrM5PSMNegSOHsFUL
mQiCy87cnzvO0m+4XLdjOdzbMkS4rtVewfpZsCLF7THJcVoRBPkGv5PQhoBeh6jE48NR1P/DTTaK
0Wq2SWVdnIAfxuI5Au8YTWmJsapQD/8PIt9A5wl7T+0esXGXpxBimd/DYTZdZoz3HFoY24sWEPh3
R4qkYZUR+Z0Vn9eeoEjtE4/ao1qegYD7SNk0iD/E9JkQ/ITTNrtUA2di4Z8Yx2G6arzNijfiZkay
FQjKRTzOVpnn64GbW8nNPIRcTFRDVr5QwksUlSQpcwU9/wFRtCzyJZO0sRzXWzC4zCu59alnNswZ
kmfE8TcooYjub2/FxpciNN0k43Uzvahht4UUr4p07Vzxt/PAuy9LKCuxzMm0UDL7yA8qLY37jLir
CJA82icnIlUiLx6OpStACPXWHOjeI/UWYN4rHrxMmUMTQ9fiKcLA9kHzbueDZacN/RBlO78vHo5y
7WyNV8THuQkZQ0MON7Q+I1AjlFurAH/btpr6DvMiI718wibf5geH9gGuFTxtwSVX0X+wjBz4PulJ
TvR3tnE012RbsmrNcOUjgfwp7eZ2nkhX5pe1tZ/TMmJlHXywa9oBOkd+rwUxx4kXwqEflxEWcDTH
fVcwsSZ6OYQKjm3pol2sfTTIE+crKFxebOHkvb2HIb2JwzHfrEvJRbf/QRTqZrygXG3GK2/9pvOV
xWbtJaokJsQvMD3/WBCHDAgD/ksTyOYuqo1zTrTjFJ0fMaMCKGxi7ltXD4pmT325gAmxtMDEMSjo
UCV08HQcKaZ0OQ/EMLi5GLNI7NnVZLLCvLweVwvO0tfAlz01zsr/S6xZ/DKjJIpIYydkpolibYCF
osOyLEV2CG+6tSDtIb3G58MNMpnfrVvfhVBFYzb7ykmBTmfMUx0mL+qf6ultPYFPwHXSGsn5Em1A
VJAW69ODiXkNdRWESdgnGip3epmKocnTo8Pb/NtiWdccFUzXfd0H/dsSOBAVJiasjIPzepgfKH6K
MhzqID7WmndKfODlEEmeoQGLE3OQzJ92SIzReY0t12huwzNrpstiTwxiyaHi5UK0J0FB+lghdLwI
8UT0t6fWzaeayExUFVMb4ekixTTgTL8bCyCi1BMrJtwB+IPJ8qJ68RROlmfcnIaiz2ZipcRWjTuz
2EYeFjxeIUux1Xd5K+KmEkuLX7hCPxv/j3VBjLLN0etvr+zFWegNjZgvlWCTmUPFvUiSCfFc3ugf
x4tzgkE+DaAAL6Himvb2PLHcNqa/EcE4a8h7R9EATuAAQL94wppJazHf7oLpslhSOyvnERvumqff
L2G9m/HLALaTwhBuzm2R2Sx1WN0Y4vMH0HP+Y2HhU7xImb1l+5WN02C4VpfTWCPq8ItcMkAIMKSd
i7JrD6tO6zNW2YdMRnQMs+mg0HQKP5mzYkmEGowPVRnPKIGi8l9ndcL9fGgx7Yh4/W+t+vm0SoH3
eaG0K7Ml5/65zoQQ4g4TBmV5ooCBlleJnALryakB5RzXNZeBfv/5hqSZN22Vmhnl80TbGjT7S78H
vEjsT4Aex1jBsVpw+POim+xcTlPJmmBfBjHWH0U4rqnk4MqUnEFHbK6ZZ/RRZFEjpewKgAjZb8wJ
IEh+1djv9T7tMRBZ5J5JFmSs1apq0roMXFtak5VVCi0G7wyLTdyUM56JlkLUy1MOmniSA38A92dO
t0UGF2bs0gGH4ZkfKat5tWLKqtymnuNtD7Ra/mKNTGDJ0iKSZGz+Ayh7/ulImuV1DQf6hlI6S2ub
b7n6KPmN5zYGqfaAF1WWCOcdYhSieAuIuIxFGrmk49q6KQHcXmDAeyUsodY2K+DMmXnexPdgWo76
NlDYBMcypO28WzUuzkq8Z28voe8s5I5ZeC/pisLOmW8gJKbW/cOV43mndfe16tXTAoNDerL37S8A
2CeP5hxjXvuvtvRjNVfC8twxD1L1EakoghzmPlJX9U4ify4C3iuYEbLdhwD9+fdN3U3BNC891Rdh
0W3jYDFV3+BNbIfomUpuVsRme1/XoucGDcmHEWcmpEpnXfD1UUEP0tH0Ro9s/xvls7A0iUcrlSUM
CArWWEKpBwnbbVOx5+l0/0iAW5vXBvT1ehEbfyaG+Ht8Wt7SIvkXFDl057OoK2/dw2KXuCgtmVF8
KzbV7SoYA2Url0kz+S6JUrszhzQNVx0vKlauGmUbbCCopV/5h5jZQbjNyqUNP/mQ6LGF1qtWmPHP
7QeSMM1f2BWc6zumXp4J6dZ1t9OC1M76kc8AIaOqLbmm9HWr/iqlJmtmRtlyZ2uBBat8OZrZ8fBJ
7mKPG1amM7QcTvbQmQcbZL3jVtiZZ3YopktJnSXovAMFUybgpEjuojPhEj2LS7tIPYuWlftec7Ua
ZQruw9LfPTMIkSQiZrQaUOcAY4TG+C8MKf5rPsxJaTzc7iCacjgLfNOE3tc7aD5oQPKQ4gxAFD3B
/oM0hy9JwkhFiR73Po0YaCOmDVubHhas2EMk8Caa7T9FF7v4F73Faed5sD1wFPVd3qlLMcZO5RUg
AV2wGfMDU3DiNCTZtWHAMXQjHro+mWdEV/Xpj/qFyqPkt1ixjVIIoyxKaf5VIv8MHSbLpTjcZc9C
D5eJ9J/EI9jkqZNnjWsyRBt/iwc+BNwb6JkdnRLbeI86T+Qapdo2xzv9PY9w5C4DU//h4OyLbdmb
/CodU8oLf7i/ELZBrQIghJi79BiOz63g68mK/iTmOipLYhBz4S0CC5nsqvB0hV21faAzDnHR49Ie
om3jUSWMh+jV4/IJX1QI3cHldirH4aM5Ls5wRajmnUzhBq9ifUG7BO2H1iwfiYV7f4yy9D/DlKIi
qAAsAJCkTvkAd6+N3VW8MIDRWA+xs67nIB3m+W7xTxRVFbpRkcfG//HepPtaDDLSDPYxkkGjwO8O
uXmvWpaDKMsfv3F+eSz2fXhsE6KUhO4AKZnxSXJQr2YtP0rnHlqb5EpYOKpNpxcRi/3WRDLFjDwB
anueIeKHayGAZi2CrgrPajfspI8RNbFbYm0R/lAGGkFqiOGSEu2ofSyu+FFpideZ/eN94Ui6yvXG
R5yqRmaLUBPnV4k3RX0CFunY1w5Qr+NlFMAadg6B16oL5XFSUCClioUHlIEk3OKlW0Xn0MfvO+UT
247iqoQqEXv6HhIJn+TUgIMM+B4jU00+uypUubAXZCjGKfKFqPZqfBJFh1ufnmhzkNA0u9qFOlS3
gzOCopa9jNefqne07Z82Uzm3kqrNoej9/dzJo1tNoCdbI3LWku95CtivAdO+HwhRQEM6jAnMwmJB
BPV4HyP3i6XVIJ39rgE+QXVTVFxJYBDm70TeHTpvx/S4YA1MRBVKcXtSKNqilN9I9nvfqYgBV9y7
LQg4mU0WdrVRFUbXWhNd/udbg5Z8fUB75Ee6RCagcUk6Ixat0qu+4XlljJ50YGJVbOvmch0e2a3H
iUEA1mVmA19/FFyWXueBFDQRYYlwVttGxUive/9N7r1Grrp1mow4N7ttkICbbBgY/G4e3c7yzj0k
e3Ymc3ebMorG4ot+gTRd3Q2GfSKeIKkDF83XU8OUi6K6MWDvSHqpXVg/2hL3hFtq4/zGGbWjs5ev
b/CwJxYqkuVauZMPi5D5DgeuHyReewP2AFgFGEnDJJdmK6k6EahFmm2Yr8bcP/bDsBey09Yl0URp
rx4UsR52Qj6NDg25xS0bxhZjhLeCTugQDRaRYcWk3MsX3rGobmWNYUBf7lVC1BI0UjN6zw+gIhn+
qOXJWd0/Tef+HUTlR2pUjfTjR4huUYM4Ufc7v/o0LNkkx5qY/KPbkk5Ym30SP4StFjt5xCTKEZqf
PoPom5gyHTOHO1kg72jggwX7FKBh98XlEhl/4JZUKdllzcWbpM8Cydprwff9wqgAwChxGLJUAtV6
wmvSxR8Wo042mYuXIfYBccM34KctcENsXUVkg+MJrDmhLNFNvx7AEOpPi1eiTPmavm5YsTTWgbn9
leleDdeoDgXpZWxsHBa2aaNtWZ0ZhnkEa8eqWY6C8awAlsffrE4mITcu2XbQ3AoY9OVC06/UI1f/
RqkmGuQ6rT6s1PnW8iEg0k2lrfWeICm4RyqnJaOuVhkzBA9XKl+5xr+P1ZM3iqyDGv9yvaE0OIIH
9djQl4AxV5HTpHBgJ6kXfP3/iM1R5JRGpCB8cvg3T0Ushgzr0oSWd5inoOa17chHGvIZNBzttCTf
5ni4npTAT6s1RU4LAJCKGLf1Iztc8AEJT7Y6Y3A2aDlOA81Ddg3wP/IHP0NHLJKxPRJBYnP9kXSb
k+/ddiUh3qHAAHrGf47vY4KeKfVxPkzQ1gTU41gsMYfm/pVMvoVQxyllDtfiXm3I8PnMQ6RHztiV
6AKC+VeSRdGdHPHth5loSJ/eN2QrkS+KxW4+rLnF8duY9CtDYCrNj/cfZ9XTyFpuI2rYCiwe3YDy
r9ntZVLQuol7Dfqzx3+P+cooVCsnTF1LzKdZOQmEnP8oFELLqJZWiPFwRtVVkmf1TDD1Dm5Flvxy
/0Mmkaiua+bu/8bKfs6YvYEL2wzcCVivJaanPSKj6zcd8cGH0++bHeMZDrVBSAinBc2UyCLfiZgP
IblvrwZPAnh+sFvft9/adF1M3wKmjc4c3Gp2YeHMYvM9IJ6FO9SIx9ZLEXYLNp4zP014uFWV4Cpl
0nMCExDGRdvKF4H3mrIPQtL+kLT2HwARvHNZ4+wD3BzgCc6nGG6c7zZTJXUIgj3Rx7xYKZ20Sx9b
CF9/nykJhQwKehROZErLT6Xn4CI7H2FtTyGLsO/T3UkNqWHbfdIGpU/b/Lxy1X0zf/h26x+h0fzy
lDm2QQIrfDEzfb+Eq+PyskU0NZ60Kdavbylx+bFPv7Jy950z9n4g+BRvQJtkwJyKOpNwvMURslz3
YN33EYRjOZVfIp6M9g6SYZxJdRVkvjfJUfQI1MB7sHavyfGfWXOFy88wAvfcoUWAhQpcYaglpPUE
wbJgubkn8ZEj09MjO51N2gNQJ1r0UJxDdtDhovBb0RMFRSuTcPbcXY/AqaWPBqDa26I9Iu/mIMcg
KDI78czF/NfSwoc3ECRiH7s1yS8C6s8f0RKw7NrbI+d/SuPBWOmERGKoRi7R1vESKSGcAAwrubpa
LFOYeszZzgNaqFDX8Us2wVdc4T7jYiOJNhG1+KxbvvZJje6mEAg2HpSJfY6CXaOwEaeq2FrUX8Um
i0PDGp+u7b64dt2y+fvZL6C2wTazhVQKtdLtTshxjD4mRFdh2YHxUBr19chn5RbkehPQ1ARs33Vi
2tjJ7Az6K+jqIeMBax/tCRstm+YRmWAmODrtEdDXIt5MSeDzQoJJcvKpIjZB12R6XjbWIAtrOKod
aKlBiIe8GvTFrjHcL9nfT8xB6V3kCQ9dD5N1oleouF160n4yV5IF+L0ZgTdgIT39c1WKiK7otvOO
DqTe2cUR9v+8S04yYgv3XQQAstKlktd5oQBwtmDNULrPOyiIRuV/jzwFZvkEED9RO0pAsF8rLmSw
BZP31IYjXbhuQJnTdEygoM5G5Rs9hglSwZwTzXUTnuQklfMiQZTkxKC3VOCifXioMO8BzDBSUlSa
7JWRYy1Zf7ez3F7FDTcj5kkRJe+Gtrjcl3bepJJA04+wnocN0nA05ZDZWTAIFLfnbNZYi6m+ByY4
/wTjtW9tbgajLOhVKpgtjpu5jWJkmxWTZjF4ZIRX3COXD+gVdRwSPnSPsEtmk4J+c0HCTn38lH4r
GSDFQL8w6X2smRqVNUunlUqc8ugAmcEKZUhdaWBV6/+0DfpgUxPww+5Yo1To5npZOsLaHkg0WMVU
elkqTMN2yxJ6A9Pv6gHdtVcMHi42+uj3/G6+QzOrlobKCdPbSWTSjODvOdUUiggFwifUzzqx+hsk
kqLmLdrw4kUfvh/y2IuG2jv+nS1DzW3WHudXsfZ2nKJ9Fnn036r49QLmAqnA3NYgbxgj+P1IOvO2
HFe4E+xCqCVQtTssdgYp1XojaSzFLoQSoluNBmvhPOjt3ALYlrorlPcxaP+eAdCW8u4mqO+6HSfl
BfCmA9PqNFwOxZgCkWZ9oJRWn53N6yWO0oF2lOiexg/dAfkHaFmJ6pEGQm7dGwDTbNV7qJI8NZMw
Bym2OsWEWi/uApVROJYIxkO+f0sJXy236FEpeoXAZ5sjmbIRmC+nZdWsiEZ9+r1ZKK+t62lc6Gnd
zxlOVEaVSLyRUi20bTr6M1T/EimI6t6/pGowUMw4WIO9kUqqdvPG/uPTdMPGFxi8+Pyxu1RkeeSu
LKv9XwoRfklgHugtJVDjMuxd0FwoaiGXTy59C4FRb/5bZFMIf7IHlSNtft751zuedLpV7sMfQZlc
MdQWURzrz3dC2RHyZfv6ImMCWI9hC/OtwqExaYMQ7ddkzm7/4ZoqessuZ5KXE12E1IirT3l7vIFS
RB/iEXyH2XIOhTgbPrNq21GeJWtfoKf+N07KucR9Gd2TmPmkUPd8aHYX8hEU8BtFYi+H0ey6DBpQ
up0/vfNcGr/aIH+4c1PdJZhv8hzqdYeKeGWY3AQ+mqberTKvmwNedM4CjaySIjUWCDUUi/k6z/1Z
YA9ffzRX+es5J4ACx9P+IJHo+HyqNxgbm4uCyxTyHQt8Ajp2ZGN7sPyudSUglOKAtHE0A/Ht0hEp
kZrEoVNRpnFplCQqHLxSK2+sYAyEZqM/affAlg08NGqFdQia4PnFYQdi+ywE3IYQeGMJ+y845OC3
3TZTW4pdsOzeN+2pff+Lk5eqtI/o6TH6kPvkdJSI68KtwB9t6aO4PY3RUAY32Oq0V6hLPTkyS9Qc
RHFVnwtqlpji9wOguIVMPs7noN+fcSmVE2cgLIYwDC//YyFM22Q7S3bClOlgRaIMGSbCsbV3yXye
njUc+jdMmf+ToLGa3UO06IAmBKTkg0sXLscwEbPEPBFPjW/TinCNQBhwZtwOdjn6PFTvrZZiunZL
iASRBhJBVlOVZaTJ9T/IuptnGvcq8CgTxPwL/m/dVwoI7Ov3otqh6IXearVoE+wdZPcIhTXacNOo
4l9SNa1BKwdP6mBmAEtdkBfrVe6hjYHVv3OIoldPBYnPaS/PmeyZ8vlqCNqnPFdTLTvwN1rYouTR
IbWpIlQopBpcFsB2XH5ved2MCXfZaLFxubOTArRNMDBD56KrHN0bvQO8xx+Ian6YlFsAwTeP5tZD
Efb30mIRpSIG3AJzxI768BZApyIB9QjO8+uFCt6ix57PMJ3T5GPBm/AuPuB9Bxy+/6avkAWKWGiY
y8H+XXgSk1o/tlAhCFgr+eqEXhxgkqKLaHPtg08MAy2G0a1IQAra7Szad5qR+Nn/tFDw3Ov7Gn9o
cIgd1XYOvdFnGFDPv+SklzZV5DHj7+tchjn01oy785SE0unSsgZtnQxpFTg+7LpDY+PWDzw0pdu7
vfwDDlOVr8O0+y/DeFfZmGhiOjCauQzNqOlvr2V5orYv7VQviDrl7j0cY2Z20nw6IjuS8ihtoe1v
ed+Nc9szFxM6w3sBM3AjSd4+0GWxqB7oJInj1AmTxl29kTPR7/oWy6YrvNjfBxdVPqgkmzh819lx
kPhBJyUvBVgW73F6U0olkEgnFWWAj55tfiDIMCjP53Bh3uj4QFlW5qd409rZNXv/eOt6w3afrh7D
XMp9cWksXQrAiKx5fQTHGXxMaIQcxKe4xqlTC6S7Sj1ZMpOTWvthOtzWFDRQU30+8lv0ekJV1tV8
KJ9fR5mYKb+qa8bFbI5V/k3l/LuIhaBmgO0T6gRXGsZtvJPCRRxDSC26CDz/nQvh0KMpiSPIHHgX
xk+FV/AI1L74uwtcGXf6aA6z2qM/M68IhT4X67AGRF8IEFCrWirMDA5QRPV0QFKesfYXt2G8Rnir
jebwJDwLd812x36WUj3kWf6So1no/NAk1BpMqvGT9HIgvPD8/WeYYr471yuKAR1lD0qJ3ll2WEGu
8pBG4by9k1PgWK/kot7nzEKQ2buppBrRD3SrHLT9UrwrytKF/KJXXmk6fVLycbgM/DZ1WKmHuxH0
hQMfDSULNfsxOKpjX5jPcsRlWI1GxYtbwQQDWGg74zX6MzuZwDE3az6nbw0touEK8ATUf68TQg2e
9AZuilf6GIq5dRsJ5MLtxyUsZsjP67IizW2Z554zZYDAsyJBhvqGbNmRh1TV5QWlJvw06v3lLHTn
OfiGEo3m0HG0Da6LhPgRUmg36xemjRlkBc5NPFHtKzV8xT4sKxLFnKEtzLZLFuQ8Z240IdR+06YU
p/eNM1Zql3reFqV9RZ3xI2vf+QfyzADmxyAdAZ/r8gSkjg7mJIC+aKYTpz5D/3ToIef5xb6ir36O
yvsaVKI/qJao0OdG+9SghA4fB+2DbO/0lv2DZvAQCaaptG+m1b7NjkOCdAodLYNZKdgzUIqmHsRR
fkJ/VRqwFPbhILU7J5Q8TC4vDeBfUekEYlTo+Mk5Bu4y4sUXe2COV51R6pSZEv+3hJ2Wvozms0Vn
559orOrCqvxllDizcSpYhbGVceD/oMYRjG3QaFvfvOSxifhARTM4sgTqqZQmtxGd8BjfiNXMiurE
9SodPU5+IfCVhNWurwxc72fKw82rAT9WQlTt95aYAtZIJiWKClPHBdrUZCbdF7IvT4Fe+xinsZhS
uomrQqK7Xz++QPfU+4h9mYJDC1gCK5hlUiVJmCNHTNntZAvD80HHIQpqcnHwki9Id8AgN+r94Ncf
adXbOkDrtttQ99Flz0Jk8CLqSkWXDeR9GB5ocWvpg3SXhuMZaq3g5peXHwQaDhIEsuLm/OLj466n
JVje2BRUMwdSlJ8o/MZB2bc1+K9hw2zXRCsLgLt0aU79ejVvvcmk+uzi+DDxj6FRNlu5/IK3bcaO
6aHVwiKtTe25TcczMsKMphYlX0P2yJfMgxumVsM41euFpa1IH3RYLAoEWlqnyY/gETxKothmHAJ+
R2cW/r08xzmD5nKdXQmr65jlj5w/EXMlhtaXUEbIpVK+s5kBi8baO7W8n8DV7ZBrnxvppwOs0AHg
Uhz1Hs+O/4EwcoG4fd9EkDkE6aLxJ2vOgQPBx5wIsPiEuwkQAyEspMl8rIesPV2Q79q1kkl5RYpC
aWyexqlHrb8DC3tt9zZEVPFUudt57pQGL6Yznb/JXzp21/iisKrF3dNCv0Hw25kUCZGN8fECp+EU
bMm4UXI9PO5n5ZrXqqqBcxY+TiigJ9twD5FUqRTCIketDJnU7DlSskHO9FTwTjVzFRcBdDeh80bX
nE7EkYHkJiIUZ93JbqgJg/F/eExnULDfvqPqtm2WNcxey2niLcoavzvsCmBD7uSgmX4cpw9nVEhH
vTKwNP14QNnbjfRMMi7IJIc3nMaoTOu6ugfBStdpnftEN4ga0u6WehrkKVHEN5X7BYGQx+tcCy3V
qxV2nIbh5oza4Ng5Qz5tfSq2Zqk5qQAdEbZEhKEwd2qobvVLtF1w2HCZmufMMKegze7N4JRXiLZn
nW9Vvd0VtZzV5jOiIFEjvWlWxSiByfMhpiMLDarYiu1Cc2JFEBLKDGaMp7bSM9++flHHYgYokIpk
7SizrKt7aqjENBQ7RM/xDbZBERH0uN6fEo2eRlDbZQnWytNemDHssoCLcJlxVKkb8FLGKEi3NODh
ePfv3b53HVJKTV9Tq+mSRVpTai9cHBVJzlvKX9XkNFlhQYR0WsU10IYjJMDFPbbRabz44NGZ2nCD
8E2xaJtlIdECdbj8n6G7XQXvrfspq4BWe+tF1jtEoXiGTjrLcp+KiGFMT9pHAibz8mwNrphuyT6w
+ekBDBhFj0xOqY4IRZcQto2LkWscxigFkc7AeIUpGmJBaSJEVAYO4HlNTB3cUPU2ri051RD03Kjv
rkrcq6w5hC2cvk3ZJ0vEqBKxYJ9zVXpD/vfhDeTK4R7gtnCB+Kau/g9xWro78MjGkLgunGp0DTFe
UaRNp+/1QIT0wvf+jznmOJhAZem6vq29usMQNnyYZvXhmLZxE56o5mtnIhqgLPC9Qs3HwuNPkpV4
KY/gsIdsUhvg0cVJKzL4SCw5vPHGkun/YUul5L/pb9oYLxj/8C063/qCdMnDntcGH6klxHlS4ip3
ynMPhoyQakBH7S1pK6Uoe4InKJ1Ldvs2NqojcyB9PFerEXmDhGiDC+gG6cgH24Tc1eC3Q7ArFBEH
MJw/vCJjRHH4AjpLkh7wyxGvGNfe+btJV5Nrwogjhg5Sb5Pkn9KZUisNaUpsXNwTBdpCqw7a23rC
OYTFTTjs+RtUsCt2lRmQMjPH8M+Z+75GZch3OjRlp2VTx5/vAKdfJ4NerbnKbu5qpsKcBeiILNTU
kKe0RCg3m7oSy9H8jAPsCYPH0pswn0aArGWcjP8faN7OaDN28bAkzdWOGtuntk3QToWuzJrYhYX5
DzaXhJPntaEVME6tcmHF5Uf8m0JDSrWYotG555iZLdd+75Y2ddxOlosO7pC19vFqDlpQoA89fO36
w7MokixUIbbs0VB5BwoVsU5p24OprdT1109131+tTZGLHLiEw59xcJA1aas7WilvUDmjJ8vyKAMS
1dmglWvBLpCF0iixhCSV1nbc36UlmV8SOGPhTwja08BeJkEV8iI/Ac7m0j+8F6ND0BJfmR/TQxBx
7HXAph/tgb4uN1xw6yHbFPN/2ZQMNFRBdhtHOcQEXplrX64T3hxJxmAGc+AE50IqZHfO/ZDjpy/U
KCNr+HLELp49uUT2D7hOt9yzIHHlhb6rywAqM4UjmKdb6VIOghLPQYUcoyFiQbq+Tc+BswSNDwHz
0g0SinIrCnAg7y8vFbPSaw4PNY9LwGfgvS8wruaRj+lFSOxdElGtnoiZpM792tJmIotGJqjBEakj
sI5+vHr+5VKwGKZl08nJ8rPZ2/Wbu/F3pzVWOQ1ZkA3cA3q77+FmIv6H1sejkESJMG2CCUHI1h01
illpnSUJqh9uVPgT0WLL3nofBCTZNZnkWm0l89OazPLgr0h/IVctyBZtXGWoIkJ41QOdqJzC6btU
FEFbAMcyo9CLobURik3VSPUoaXTXCBw8m+nbla1Cbdo5QHYquRKbTX7bMLdIDtvJYsMZynzgOkrZ
aFsWIWAqGVg2MeXACWg/CL0QUrFih+c9p2hySwaG0tgYJgJIuG6aQsWLbJeUyZuwe8zxBrntfgIw
CuviDd6IytLkqyjtdmZ/j/YAdLdbEjxqpLhuGhzjZthqoWgg9/S0t8zARRvGtD5ipMAbRuDkDqMA
F6MDEefVnzNg2SvjWJkGzn0ISEcFL6aZ+wJKlP/ZBy7wg2o4+dEUOqT3Bvvt6ujYk5OoLJPwjcZE
xy7c6UNwP8ycgzkpf+PlrtAx1eVN2VSMvaCtUqEwaAbpu8p3BOX7LUkOHGuMg4q+E6hPVsnpITvx
DRF/kCFgP7T8sxlXzBY7l+XbFRnCr5XQdUoSUwBATxDGYq8U1p+2sJi3OQozPrFD4J1bpgyHC3Fe
cmCxTVCztYWVlc3rB3BUJbsnRQQAuVxE+eq+5s6EUA0cITYPw4p8GcYd37n9S2jqp2yAR2rlPp8v
KwU23VXco/Vg4AIs5NJA/D5CtJLeEzT336gKmP6Xkw6NQmGtl5OAmj23/uOvWca6fESLPjjpC7bq
PqHgzT3i2s5B1CAq6IE5YpO7xui8bsRogjJ8MUqpfgXiujp2JpwWRc390ENwes9yrXc4enzyLT41
MyeeQLg/Up+lBaHYeEAgk36GD92w00bV3ijXA0Urv/m4Fbchd0gVyD6qsYmWSOhOm5H834kXGBMZ
2MksnJW9149ABKQAolS5ALBRo5THwyUsCFr4PPQkKwySi5XiaWGiR+maE7m9JUl5MF8bjAlDgIwW
8jA/jNytUQHdmnTLh1+T7Mavb9zeveT2HYZbNcM/6VZSFZj9l3V5UkOg9sk+JCvRiModKlRRKesp
wQxK41Y0rYjYaMKBzS0dFPg2Ff4QKhwu2XBXcWA2WtCslOn+8x+Buigml9DFN+iwbYvo/qMiircz
V+lZX+LpdF0YcDrxpcvreHjMxkGXylW7khMdzZ7OdYETK024mikAusRdB2GK7b4VINkPnDGaD3f0
0Qf9DCILn+fVxVJYDlOwRWOTy/jM8bowsLFmvSkOd1trJM/ZSP+wTI35gpBb1YH8ISJPewIohtsd
tWc/VU+I/Lqf1M3aCVOI9HJFDJd0/EilkGXaXkZLKwxzIRDF1BoCA0rfxbA6N8rnQbz9HnPB/8Bh
+tgHX74f7EtEoRp4UE7hBfKfGdrnABQN7covrSKE6PCEVmLrdpqS4svEjWav9XBuLGCeaDwKRI7L
GoOCkDvBXP1NqXe3vL8fwBD5vFvvoYS7BNMecvjxZgXq0QjZbzNz8389zS7qC7e/aqiu8txoSifr
40xMxccTfWB6nXB+GYm+9QKfyyoyuF/0flRshZHslRf03FbjvYn92/a5ycK2BTIYHakNShKWvi02
jHHAh4gjtoeU0ckvY0WckHHItoJk2XoxOneA4RqA4+fGuWx6HE9L5mCCWVDOSVVR44jkB36f7nSP
INKulsm6WEar8GX3lPoHoE5unErlZWOLRi8jmQTO/jOLdIK39HDoimw3g18LRWRqbEQU7zQTcyQh
0yX7uDvGkUERyTG6lwrvpm3+Wp1QW4mGSjrfXI2Y3FHOrmJTyyNVW4Dmh6ASIlUKO0Wh4AQ1Frvz
MrvMKKG75YB/H0CqtbaTnHVTG2oXSQ4IGGbk8nw5XfBFIDHc+tCPkVb2+rcFEVzeRdsceo0RHJZS
9BH4oulowbvy9bwMgQTFmUf5mvfdtL+UV2dkSGOFzChBT4s28mpI/trvpzPNkSmTuC61VR83sKuQ
Qvj7CwyO2iTKcGzNRCms8O6CZqm+CQM1f8sDoNyZAIplOeWmjn1fw+wcc++CdIpvnzD2tXGQDkfv
iJaFPL2vS/80ZcyRA/WgIQmxTagVtH1QqbX+/TYG5q2ldUAJA76G3by5/vAexV2tZcMJKVAJUn05
6LoGTOOgpf6yDtecpaIwp5ja8lJ+/uqT9i/d+ruGxhasB/i1XLIMNx2alSqrjtJAfLPaodXh8EjV
8c1TnWn/EYpcicaKl9UA2ATU7w5lwEiZYX8wDFVYY22gUWb0Oa++DL96kuViIFAyK+8/KWlDML0g
oFstew4vbH3jTM+JQ7YMocHVe5SL5AqWo7NlU41g7pbUIRXGUsoax7gqV6DGAdTL8ta/M66K2+EO
6CfEN3E9pGfRnWUGgJJqQPWeyVd53hBs2afn1lp9WhzlDJVE4zwZxzDCijPKxhhLSUktCMJ0GVU+
JM/nEgsjvN054yWB9e8mYUMalmJT7aKklEzNMcOHL5ONHIDtm8Okko3See1PgnJulu/2B7oyLymA
bMP4R2cgsR6TZ4zmQBxOMuw7kYzgHAKUGj2xkPdGxkpYQ+kT+TK5qNibZECRj3L6A0pJ5wfeKJ59
u4OP5C7elDOoMftdqaZG2PeWtAVG1qg1Mzg2K6wbUnTGHz6m3nV4dvagd+6xGJU0u1pGZPSjeKnD
7htuilWyWonnnvuzaZ5IJU80IfyYk/g0/PKGoHRijyD3X90u1Z0Gsy4dGCVw6+jBkR2kxZT1r9UN
txI5ZAVYDErbsL8q+oeHB7JTaVJjUekeqJkAfQldOQHFSkoLxB48X6Cv3GwjeqZo06dg6JOMQP03
a0GIbh56NZPyu3w74z3VmPQ8dO3L6+YEPImtQqL9m3SkQouqnORi0PC+cdittf5hLT3ODMAZEcc9
D+GHDQtj7eRlf3ucimA5WHVztvSChQpc5eAsRSKWVHeQplneOo7meECFKEa5rsyBMWxeUNvgCcJp
Qy1dw0cJrEugDStGrPSlA/srzkqcRKVHTSoYAMlSUVI2KaujmQOxp1lSjKrDUfKLxBbt/M45gtt5
6KP1Te8/NjW0YzTVFqF2wGKdZ7TENRM17Pmyk6AhosfIYFEBvFZMMRr4MnOl5nuMzJDPHXTmMRbt
C4wNjqbNAm2ZQuCuqXgqA7eINrdclzJ9LToNkrVtBQeOABVU9+ssurmxa8nzlkOjoc36Ma0f1dnN
9wEKlVKbHzvES/QbBK2Glu/JmiEF/QC0kgyvVD/Zbg6DX2iwf6vFEP375aYe6N6yikuBMAOZ6ne/
t763FCPA5/rcntHoiXtVqS3KI3PHE9Alarsafu6RVrWhcUVRgKPtEhl8oNOWXG3TIUUONUoLk5T/
eBDlW5xz1D1X9qbefD8EBae77xEjkqGumEzKdgAAac0O2LGjbaKf0JtUNdKfi+X8ySFivJPxgItc
+S/Qpn9F1TsExqZDvCbEAeFJsRDvSzlqq6IQoqWiGejFZZpdrvwAehqzlwI/Ls+mHw0vXYT7heUY
LNvZgF6JnScEC9dzSP+iG4ZQQ9DCAp2Y7eNlipN9+hYMYObBdaP++WcdmlYFXRqykXNmfg3/ykVy
4jbJ6bz5yB8q4M/cc5U3rGtR4AQHamhgCJ9sgtj97StQBz2LnryWt1FoT2XWV0KHPfSkF/m22TqS
ND+ohJkME64usyhgVhVSJSY8CVKiWRxTmq4Gg9B8UPv5ccEuQGSYl34vGeZMkMPQBCqeqW6GI9NF
jJJAaFF99Y8VRozfjg/0fnumKaHLwBCYUmykdSetRA91gBWslMR1csljmc1c3ii5v/RzuHPvT77V
ZS4rYO7dKP3Suupp+EpCEpNOT0a67LAshtFEWanr1Jk0tmCoLsZfSfAJJlDpu7K0m3suFya0Wvyk
UjQggD6Oa1LR/2tEbSDAEwCL/sgqDUUpoM8XUWG0hfTZYi5hGPSJ7a2BMcrmEcYwgv4Qq4HaeWc6
VwTI9lHvQD2LcDL8buSjc5frmXc8ylSLxMEhbnq29loZ0XC59b9PTDbRcGadqeGklGSEr3dfjaGy
wySetpdYYWDI4OT//FIobmIR/ZTJtWpznazqDh8Te1OBU0LDduTSuLvF48Ek8gxFmKLs4Q2hCTDp
rUBfUcBkvjrLEyoIg2ybkh5lir5oUzsjyvYXP6S3LqLlCNkT4MH0AlJ+4kaAsdfCgvN65iRyoECz
qSujwlP2Me0twxOwgst1b2NJZ98aiKiq/LpipVThVOJk27kj1oQCbQ33vM2SEQ/LT3ITopuKiXjJ
z1zF7CBMrGWB7vQwJM3TZpinoPDlMchqI6Cmq4Z0rdYSBPJ4aDRMjnt0VJCnkQLnk/Byi5rB4VVN
HUyM/fOgWbukmWsb0RPDBPCR/qNAc4c0+mEAX7z1Md1TAk2dDrdPWY9BzdfpfmnYfQ0nhtCBzgQP
9McIjv5Og76aWNdek59hsHeRdNMvkm+1OQLreWX10TXcPP9psXVUP1eh75y9o1mTOvgPzB24KW5k
xJMgUW0TEfXLAFUY/2NARpEVrjJnuZMdc8Sw9jVcaD0OW644FnQY+6JrVG6rskQ1arh2/joGPPtN
OimhDXRhSj2IcBYPQD/72pTg/tL8pQkELGfRhkpFZq/Jgq3IW+aRtjgUgEphi3dmC6rRFPkyncIY
pwd4XC561pfqI4a6bK6p8GOg3bzY9yP91BSxq8vh0rbeJFO2NswrDMCo1wIDwuDpto+0uyv4uX98
VY86RbLX4WC8oEWBMai+V1ETCgA5pOWRbVeDKyXPzAy8Y12RlDJLsrgvuXlYWLS/y2J9ww3JYxDJ
4PG6J4LtzFDwEehjv1Nrs+JCPR7wm8wwsoyHjtG1/IjCG8fBMWlmaArnOkOKastP9cfz1n19t6f7
DOdgOBJChNVO37rXO4vw5LqhxqHtzDAwasSo6SNdYyNJMObLSTJkpOauzGlLAdItWUse6VKKj4vO
zKRycG1gtH1tggntg6pOwGiFB1i1xVE+KcxHabN4ikCS5L8hTmX7OCln/rX9xKPoZDtX0tLM82IV
S+cq9p6Bm0r4sfFH3M8CU/3RvnkGQzstS8pBKiEt3pJrdQ1k4KWnPqPa+12dqDN7P1HSxfry81bP
YaAeYDYFlIP08VC6/MOl8N0Sa/J2bg4NsSkRoPUQit0sbpOm+of0N4UyQ3EdZzGYRlikC82VM0/0
bB7iG4Vkk3c8pAEGkDNsqXv7apAm91+buW2cOthBv48lO6WWQ/ZIOSpFFXQFC6PbkHa7Qdu4Ug+d
fG6z+4IHTDPImHQC35/MpUP2+6tkL0Xhs82s8qOD5WvPJG7IZ3Civf7YfZIRblzr6aQn5qEHLV/O
222pW4znER0TH+x7yRzi0dZgF3HFg94Yrxs/aEQIhseddBMmpeSSjC1xvhpOjWK2RtGGBDvHvtLT
LHdf8hVx755HCiIbNVAFEo9fAvjXlbPYqOdAHxSjtSUggMs0LEtSAlL4Huauk6pi+aXRZBB9u8A9
4gTyA89jrCdfxPP/Me1h2qWl/bKZRdp2n/6pKsQGbCxunXy6C6uoHRK5KXVAIJeShF2OEPlZQwpV
9eLUtAER8vWxiLZd1PLcq4o5FLz8auS9tPDUaVu44XchKP1OIMPZBgrVR4/AmDTLdRyMzF4vM6rd
wVdAN3UUG1/lnvlw7bz6T653pik06bSGQqpD1oKWpZy0N6YwUvrJ+0zDeKDYaAIuHhEkBwAGDiW2
PLLxj6TWqphclTPb/bH5L8KgDrH/C2OrpRdOYWGD37lyir3/yY+5oBAB5Ng+gju7Tp6N55uZgZGC
DgUwTioY2O6ZIIAEOEcUTqiK9Bp6e5Y8f2BTFCqLZz+RQ8qZNeOGT7w3wu3fSXFHNfpGAjBNBQLd
3zIwb9cik56tdnLsPi413+w1vWgowWGOUcuxPDGVl3iL2rhl8HLDdgDRWgJlvITc+b/qPOLrqxiK
Eq64eyeeKi2EZy3q+IBk/e38fdpkQux2hQXvBgaIpPuVnoIEj9fNb5lPQyaNxk+FWEn6gFd6VyA1
W/A/yixuGjG8woqFS9cRUeXgQ5PlIGI0Eqp0Rud9NiliWPJuuZujoqQOZ9T2tuFPyTwmarEWdKq7
cMCoI1PGjVBUJIUy9idQ9/0AOk4oz2IHDgFDDz9DN5YGH70Fp5HYr3lLrwd0mikbJMX4oPUJ8BtP
MycEZ5Ka9jQWywBrCIz57D+iqxH3HcanJR3cdwW4KWaT1wrb7r/JpCdcvR37U3NrOaOIWRn+WQl3
DksvbjNcQGW4OHr2bvrDiPIyZLiv2TXHtbVSEdenZiBOMxLjHeQZCwcUN30igYgzDaBLkoDIHofd
TnoK7McZkJ4RCnHMToBHJ0NLxMGtPlxXEEtio9BbLD+IHW3iozjLGSLCphH6MfmVEkP8uJRK2jkN
NEZtUbMQBsU7t1DnxF3cjjqto2KeWe//fpshig8vK9gRgTdSUzzB/X0GMY7wkWrGkpAsx4JIBypV
AvGL7HRx1obebEo1RkSsPcUMNI4j37qyU3Fq+531BtPb0mglmCioqkBq5T2RexBotWiFZ/JfUYl7
Arjb8F5olEEE6TNjN21wDgMuw8BHyMH2uexxW8NDyZEso/FsJEKi2LaHibpFz5/CWD2lvfUl8GQm
0hh22nNfuSWezpRk0mjWDlrL75vghwgj5L/ma6Kd7MtXc1Jjl53It8N5A0P4PYaig5lHeAREWmgh
11MfcpDJ6WheM/2LnsnZ3tWIAaYbFRnkkgQRbo+7WvEevoVy+iI/fg66mmWTleZA7xbeiyKQPs45
kb1XIquz0nQcHjjNQYIC7nqXSmpuYwNZryDExJxqnThWZntb9kzHNJEJDec2+9cqDZiMQjgVxVQC
lH2CdFlzQuN5oTLx84X9AJ0pegF5cwZoXj3expapTvqgs/evsnILYDs+LDX+ZXvvRoxpTXK+6xk/
FpliqKja4A1KjL7VdwG/pW9xKy1ObG0wJ0KSFv7RAzEy2fvWwRR3R9yAzQye5kyMGxgwy+MsbIGS
SZZ1VKcFyQKBxQpikPygq+adHoqcvuszVD37ZyR5mokKx6y5h1iyZG6VfOR0bwUwZKPvb0pvgd8W
TsRLUODqpAha7Hh47dEtwJ2DxNER3ZVHq3PtxYKcxb/QtntPHe3Cf4fa8thUass1T7j6Z2UempF6
/qh7YcC6nc/rdkkRnPY0lSq3Ru+bMxCwfZVNWTypPAoy8zlT5U+sh/IDAbtoL56yEeljeqH697Ma
97pbuJyIYcqjO9Q/NxzQYEGKpHd4wQZ7ev2YtsK4zaYobPcsw2bbYpmRHvPjFaII18KfChMZgh7X
aqglNs/ecBYgKXv3vKgnMsneZP/e8jR362lbZWFUPIAd7l6Eg40l7Rk+buudvr24H3reuZVfSEVS
o9pT7qFir06eDJUF+imYc4FtQZpxIryF7/g6Z+SORBJRPI5c+MgZJnb571gOwxvyyT2IsGaVOo4V
Vx+tJxcAZvJH7cJ5BexkiP9Px+ZwvPQkInOZjuzlD2XsMvAfbuyihUc3kgXkA/3S8nZ9DlgNuyY4
fcvAYq1wwQGtqY81WUZjIFmvqHp/5umedCuCuO45FwLVrrxz+Dq9U/8gKR/5AWCXs7Bcccwmo7hJ
qt0X2pc2klbzyctkZaH+WOkmOkfwu3QkIDBMJdniB2la7ASw0fFekXhDRnXQXjZazkdNRD70Gd/y
WpLkL0drTIHOFljDHCDOrgzrxt2B0lQAUPCYac/YhtaUeSSf8f1wIaSZd73hC4pse7vYv+FktnSz
ddHyOoqSYQANJ9fvtmij3myQ6VPnSWPc/Wv++dsOFFec6fNzD3KRa+fsGNHRtT4WQ+GoOxmXKYJ7
hyH1Fjaw2nZAu0853gk2nI+ya5R8wUcmFoQsJWD5t2LwoeaYWAmoSW+RsYpY1PYU6q0SXMqmc30C
TzaV+uU8z4qXTBeA9St2zGTANZTmQ066HcDYDhXcyAzdW8U4bk7u1SAwqbWQ3whDUTgGOEDYtChp
HJXCTiDzfizGPsZv5y2NyJCR9aMKZKWHxI2kZdp0KKFYwDtm0Dh2sfmpO5oaY/U7D9rNy45rAQH5
KvazX6NBB3v8ck8FqI3OHME/IAaJbH3e+xIcoViRpBDCOX4wI9BQbO1SZZXNM/nhgQF5MJo76wu9
IW+2oojux+Y0A40kKISg0AtQSQO4d4j4hkD3r8nSbyQkqfttKNpYl99ahxB7+LHPGsUbakHwmnn1
5qSvxX3uiQ/Z7uFgPIK0SV412iwQ3Dhva6kwq1L6LVVLIKKpOvT57vtSthG0jmtfqc2hZ3KKW+sS
el1rV/CutdzqzuZPZP6sAvzsgB+dQ1vcduf0Em00oMo50PHKWma8ZUzchQmz9JI9jOAsXwctmJRy
7d7yzYI6Vg1lybGY+/r6K5JT8lE6mQ55j3hku+rdtSZNkr8D9Ct1J2dgBnGlLnSCeVvY8VoRbwdf
IPWC8FXr1e2E81fD3UXEoVgFbwE3riC6hTbDIPqzu1nlEhZcwBQevjtMhWsFy/PvnDVEy89byT1/
Vjn/Hh2wRaNPIE92UOj++CpN5GiSKDHJBPhY+klt88d6t4u94B19xTl/XXBAe6NgPKkUKHQo+O4P
xntDketXxmWzRRkgLb3lxWnbOTI1gb0uM8TK2Kw8LKg/1EpGs6hwGAP0eOXejYE3wbrCcdj1aRAl
0kmm8vngp1hPCY+NxaoDueuyB5PwdTEVWznXNUnWJkS3TruU6E7TQMKm3QJ4Io/ch/7cMG1EtTDD
1knppX/OSltKi4M+5xptYg/VqXuTKQ9USu1t8tNUIbWDopLudmFKXQa0YCbzVgFbuX2N59E5xTIE
Kyk50qFSDsAJ1xHkMxnMpncBTsGhbrI5LusVzsIZWWJYPxmz6kLgqsVgLjlTZhZwdqwWm2wth3Tl
oZeZcrMYXRUb6H+OVEsA0UwUc89W+ELB7LfTQVTF6dyv6MPYKX5Q6NLvwmOnfViUFwUPJNSkUTgd
G1vQy+6dz6vIWHl7KDaNw38iJLNL2duGvaN0XEKxV0RqTGo6YMoemKRIjVjXSXK/OT75/LqxVD1l
EuTLhyf/v2e20kqecPI/64zBUN8i1mbWBbZdysNyrj5/tcKeBNbt5bR/LkWr+VOwX9gD9jsjTflE
K/nQKGwpXKNVykrAwFk1ltQ9qrvWUpRj5lxWX0PGd0Ri5SLsUV9UqUB7sxwHSy83bwQD9u57ZQgB
IpBuRKYFwYVI6hZUNXzry/Yi/oE0tDiqCf/kHtxc46ojBGnLR5ZtfBcG6uTJM2njUWfx5/2lI+I4
I3ArDMxUEE5fJwUj48RYcp3KESP5d7dgY5wk6MO0QvCHn9eB0dvUWbTwkOi+Q04VRosTg6cVixgd
DlPZbMEroiRzbA7lSwcLOh0ywAJZ9A8Iks8/U3TQbSCfXJ7cB5U7dRXPGWO9JeqG3984SWuhi5TM
ob+5l6n3pWgpLdU5CPgn0NaTfCLAX6DVgiSDRA6wnLeC2hhV5r8k9drEaaFwW2aTczrD0gK8Zhyt
KdB8HqFqZCraLF1noa+8qQrzEmJ/X8HG6/mKLRZxqacjeMqz+ORcBBweyhQHJK6N0xAwiZ7EuKTS
YX0XSwGRpG3RKOAXOm8tSsUcx+helWeUIOVbdWSRLZeSDAT8+zrxLSs8gmIGpgmbZ0maPI7N+GOy
pSRTkoTMHo92zIwVo+nZC9/LZIRp3bNHUPXz68eEkZJOq2cPqa0qHct0AwHG9Sl1AWndPoAz7/2+
giUx7pQqmRQJ0s6fvNiVWc5Cb0uDLX8BD2aVtlJKVX14fqj5OaQCfRsoc/g+Ogjpg194G45rd/ie
BmeyWPRL1aYkOmdua0Nqr3TkJZmx/pKU9bFSem7AJB84j+ZDE5NRVUNu5h7e5ywPNLOSotHHLJXS
CthKjdzsDfYfTnOawgSdOMBvTJra38SEkR5V1Ou1HXI9Jc8oDYvdJqcH6Bqve9y8DyZ7KPnX+4R2
m1c++KPu17yu4zBM
`protect end_protected
