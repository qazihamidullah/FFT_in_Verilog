-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rNraDrxcQrNEdEtpKu829fSWh2bL/X6Sz5xMaGT+x+F1f0ZJpPoePZsQyjhj8KiVNJJZeGcIFC5u
A7VnC/+cDf+a1wSjmZFlFoaalAKYgkMCp9/+2aZaI+TQwWVYqcSsdm2KESJLdMFFBSCqZmQORbhZ
1CGB1fqscrdQ7t9eydY1fENKhBrcoCW+UsKoLZfyFl+doGCCGEMbA3szfWs1N/AXv2UiuxH/UNSy
gpCxPORRdMSiyzx7Bp59BQDz8hYlLO3LCQQFuNtZamMEppMkE56RyTAeoRi1cRTNf8GS9sSULkKb
uufTBB4kPnF/fyNCKIaODwK9tPPMEmlpSH+J4Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 45120)
`protect data_block
gASwabHx3C56TYKIod+NarXLmcn61QF6u73usb0KMreqqTRFz0ydzzKBUNs/MSlY6X6fkf12kMo0
jadsWl69fsFhTjdrPbc+o1aGeSWG8+LF/aJyaxFn5oAwgSWQ8BKvbuKAnZBy2L1rrYyq2Uce7adS
z+rMnNwm7qmlMe+INcbAc4mcCe9qDn50eopZtZokdONwwnR7Jf6ou4EtYHDNHbK5coiJu+rpUDxy
JVRq3o+NjVoHi/y7jTY5ydIZioeZVMUfeV3+Jf/IRdqRrCA8pWqmOVAkmPPHRiOlSrdLfyj7AShk
5y0SDP/aMA79u+jQxnO3IYPGMmjNerveWN0mpVvn392ALD0ve8VHKYOxwMjr/0UDHq/e/COInWxj
E/OnNBCcq0cb1x1eJxSHWziP9h3l9AWWfjc//p4msYtU5NAuiBWRuBNPlnES2kjlL+Kwok/Mqawn
vcRJzg9BYhe/RFRnUkjz6RBfsCKQ7brdMiyrOno9srrVjDr+x0dCmxE3N1/6vyjz5a3QzjWrso4P
b1No9ZJqnu7fx5O1PdYDP7uA2ejdkWimBIp+CNC0+v10vhzakbpBj7F+NCrFbzr7ptc4G722JGEj
2fTWQsYbx20ZR6B7SAPOWsDcTqNSSgXMMELd+rE+PnpZAhlTgNDjx0fCAlNwCQK1j+MdGpBmwqBA
tKl/LpdISSm9+nmhY8ECEW3ewtOdvi4aHlUnFkPQos6V74+fH6J/ry8GQbt7Lik3nPBZWAxBrldU
wfbvWSpgxRujYYtIcQe7fNCIDOwk1Z3QIOWblpu6py1uPOKfQulhJHVqEuziB9czcnWftAD553b8
bifP/FhtcGZ/f6fVIxoJ9xTZq6hRaZNx/EC8ah88PLI2FZxNwrKNNK1y+kdPidsdG+OlohoEJTP0
MUTJimB7JdHFy9xELHzgzuJLbczzIwcl6tksqhN7tSX3A3PsSM+M/fNaLaaEkp7i4WjEirEYEGYt
b4ZlOVBdpBINJBvFOYybdtz/ANDjd1xOpHXuPJ3Btv22/zBRsijXJ5shCwW9juc+P1fNILrbx4mc
ASoOxtoRwBuzVbinM/nkKQ0HUcNHkRjVBF/GgE/qGgmISTfA24gj1ivxrw4uqC+ntZnZSL+BeifF
KXglwv/NQr95m73YZcr8lUUk1bYRZW5XJqE07WLa1pbr+bbkMfoUEWpjjKqoM+ZNEInJ5vzbMIgw
S9WvjNuTR0T47sJj1ItUS+JxAU51gfKGmBNkS0sckHtVUoumFBLRXqouRzA/AWSwSJONgsdXNz+k
kwInMxZ6HNuDSpvMP3swme+Pcpcb9QzXNxuEncN7tzQ7AUmTBTa5+5H4+cbTt7FXDO6u14GZX5/8
XSc7v5x2XsckKxTKHqE4CsqYiR6Y1WyPaOwPXx0Ug3y+K7HS1SCFYIwFbAC1xZkXIgZ9UD92kG+O
wzP4IOD01MUQlcl1ZxHf031T5/WAqWSmdQXEReXUjJS1v9m1mx2jkQPV9dH7etiOWDwSbim1uho4
Pgpkva0Kfs+zhlz3bKd+z0pOcwtTiXaPvdJf/vGJUAvxX2YSO0eV+xqDLhSQLS7H9MSvsJLji29U
Cm1pkezLfvC4vxkzczlRFO6shDmFU1d45qoaveU1s1uu5/wpxUW8yrzPtQREMO1oVrdW90KucUcn
aEX4uacSd6bl/aBOdVFJwr4TIJr2wGgj7r2hl0pmtpJMGha4LRtu6PpithpXqE41JfDP0MVedhZr
tLbiQEN/AS8Ejcyaff6dxDz26H5tTVCqfnH70m3Q062u3UG5UMFZ4QygIiGmaAC0Bt/RPDM+JITc
ZO3a8bTftxBoJsek0WEGP3pxXd4F9FacWFr2aCmMImD7Pw2C+z/sEwdk29ADYA5W5frT85DuZlMW
xDefIGaJtmhamOpRK2dx3PJe/8iPxUVmzV8rKecIU2q+So+OkngidVUMr8m3FcWKCNmmCibVzu3N
Pz/7QzGvd98SloSdVFUNGA0SiP6IDrtrxEbZQfUT58Yt0/MITVgroiGw6QZv7WaMOYfjVSgQjxin
Nlc5VxEcywtE3q8IqHfz5AEYwrY1myWfVDdP2X+Ha8iB9UajKu1BmKcdzd5glnZJzwUBaavlzZyy
thNqA+0HWgJkZAYASTAd5uDb9vJ+P3yYIKZUUTxinvzr9QKC3GBHjbp4ykKXl0hKmgBTulrc8T/E
LNYDKLh620inS1c14nGZcbgf0HkHgSwzhBIDBoJXdGYlJR/tUooyICWwN1L8nRh4hB8N2kIBOQx4
QNxp52HrLnLp+DUHcNSXMr0CiG2mYzogPoiTrn+hRs3RoH6vVj9IhQ0ae09+5pEKSnmpERdTzHD9
UuJlx8r4CkWBiYwWMekbXRbGHpYZejaWZTjwK3P/y9EXyeHyYHwVCbQvCnBk9HruP540TPQwP8yl
i/OQtE6V7DFUrkp3Q+XYRz2l6i/q1LPdL7l7LWyJSDbXOqj40yoEoNpAj5cLFfw8sOOHDmvD/AAh
o/J7aKcz0nq9bCZBlDvdhXti5hm3SJQoV3eeGIt1VtzQUTITumE2KDn5SPHmo21lQQo4IHEgGC34
w+qA7gBaYuDHD6MHpoHMXIJM95zvPMBLYNRjXQmtNBSWQKgePHANSbiq9UQNaFPvL4P+bQc+v3Fl
gRc3O0RgOAi+EVznNMb5glfMmF8SfHMZETomAzd0pyEYT7ExQsBA/YH80RAXBI4hkXztBDYhV4Md
6x7wjlU9UWcpklIyDb5ree7DMZkz76xoZEM10OZREvGSP45Rw7jpKXRVnJSdckt0MLi/xWSFnPiL
fhQTzn6A14e8hQZU1JOI36aSJDmxwjG1MJAYThmYkty2fJUcbG8JW2vzQnH+QDZWYtc/qK6T2QDq
Md4zmR8jhyYrPmLnkdXg5K8J1yp/G+D56MIU4RHOHhV3rvM7bTFc3HwHrhANh8aed8Xuv+A5jDFi
lDpSqm8wapEVxsWimKFbzMpNWi6JtoslqzNeKWejy59LTT26hoaQm4jZLPV7DFPIDnNq1RBi5MUi
Km54z+erxkRg5WmWqiMTlJH8KOSNH7CZUxmgY4V5b0D+YxkoghWT++jPCh+aN9ZFo1pBY4OC9jxd
XrTEpeFheuGu3GN5Vojjt9JsFEE/3qw/FBN7N74RQRTRpPDhZ20sq3N59U82sP9ncGukHkU4mCfA
2cNWmmURlfTmWFaPakhjElvQXp2gJ9DKeoOCNtAZFFridj4EzeX5S7RTIxauQlNy7ZxhTerzuZxF
bH9ALB4gs32Qe4T3yCu4otS6BcrotsjZmHqDkJ8vSGi0EcxfSK5nQ2CQ6BAa0WG67gFOOt+E7TFy
Aoz3rQ+TyKmlYcrtMNfVe17UmmT+V/AqUXeTxaRZ3l4LyHrxejHg/yj68BYgV+l9QpL5LRGLe5Yx
3136dJtXzzRPb4SdmCPnZ4QCyqP5Dua3KTlJ7nzJVo91prG2gOlGh4CztVqhBrEx2E5Ud5MCzIkF
j8cIrJz6VFsySYvGycKpVl+l/iWZ+eMjnUqX4y/g3CvxJZXxyli5x65vZ6M+gc2JXBhVIMjIm3pP
ALIYzh1XHc1CQ8gTBoVQM4N5EbWYHigd7l0n1QhAGT/JBymQ/kbEdLNxgnFcOgae1LhwdqfWiXw3
KUPuL6ks8NVRi/6aXaN5OGfb8JdYxOgv/rlc+BqB+kqrrgqtQqwA10KeTtBHRlPUpfOdpHJ6xAe1
2x/F4X4OBp8Y4RZhQWmtyvAkihw3J1nH5qHdVDKQ4FphXFYG8TYLx62TxjA6h4SqSoFRjcni0QRe
9siauB2jWGw11ToL4L0GVVmM2hFz/CFWgpVS3grvUJAlObroBiEGTuxPnVS8vGmv35GhzP+wqlZ/
6blFsDq752aepsG0vLYzlq3vEjdArInbQvkitpgtFDFYA4A5r6Lfh8nA5WM/xl+HEF0kYhZr3SK8
6ORqscsf7OmM7uqA8R27PYcgjedyheR/CutxLd3tmiaf+yByfRK/hLfyiAqiWw+KDEr24YtV2+8S
B2gd//HavmNY3aOGqDfAmhMEw0ReWoz9vjl8YKU9JECNf1ktHhIoCjHZTzjuLL4DJKG9Zicvj/HJ
h47Fe7KaunvHPTNjhses6FvVCgqqpixgN4uAth3KdHieZonlTtt/+Tusnq4LyuW+0OQmaC0rnF7B
VremMdksL3HCm7mRkoscvpP2kbIeZTaKJO++8CdLHY4ger600/yXegouJeGpq4NZADskjYUJdwoq
yrVgat/KtyHAVNEcrUKIOrIf6H28Pdwju6tBbv5Y/YvsHrfuw9LHraZ/RuKGV0Mce4JRLP26PaLa
+Hoxl/q0YXBPRL+Pl6Nd/nex3iAFVF2XqgWK98E7MjKCehe0qNoMegUsg6/pG7b+mrkZCbFXtIV6
5cm99JkPwIQuwaWmH9iz2TAlBGmiSLVM08+/IpOnHhyP0JDZxjqr6UoYcGaPK7oYnW4IXfVOxg9U
RmaVgK16oD7lG/GetwjbsC/DW41eB2ZH/UTON94CUoZy73LxWagpxjQDTmRfRMSivapRn14+ySdd
FZNWLNC4RuvXQRBFfvxwbV4MJL1qaJSrHbsRAVuLOrFFBnBlBFYX4fu6vatjG8grzzlkNmNQMHXZ
I/5It76K5enI9iEgP1opebfyc/ooTmgQM6ial+AjNSC1QbbEFmOQjcFeBt+5vfgCW9tjFK0VXm3S
OXMcNkhodaySqIA6nXq2l7pLKQJvjwnv445DL81mhoH1oi4xZ5n2b47LsY8QfaD+3/pumciQO6B2
JNwVb8q/PX6kE+zgCf/Y1iy46DBQUC2/1h1RaCNOmxOkzTyR5vm+BYfyadhlcBe+ISyN1MsvgKgV
0OLt6++vMuo8RXTaqMkpebbgL4TQ2qQi2ZZqd0/M+Ci5veSQWgJKuhTmoz4YHDmtRzPIUCQQ8CH3
YvpAC7HVyrWcQAuamh1qw1mosrb0uwbYnE+vhCStwah4gYGANGlJcdEesne2Ti8q1I5MifYJ4Jtq
HH1qoUogNNWUxxK1XOthX3MiPiicbSGkcDbC5CGDESkezg0iU+tv9yzReKjkN8u6NLMTdF2RjX5L
GI1sVHuibnYxSFN0jKFtNnGaieNaKaiEiCA8GGh/HIkwxKtRyI+UGcxfOv5Qb9n5rzJM6A6wgUKh
nAgLbsTxKpAgaC/15P/6JAS4qwHhiiGRcHAoPUdte3v2XyUqna5wCxuW+2VGmKvcafMOOY7RFMX8
5Nt2QOP8u8beYRw6xr0qoSVKTvCtJF49rEUTGZx2DE7mTEGamahQXEJHcFXpVHHttYkRYf2Y5o/C
ONsU7oFXNp1xgnOqTK/WP0KrbDIz/0InADg9Pud9qQtiQkv6IQK5s8881UVTOmjWEl53E8Jr92T8
2LG7AT/Jq/icIPhlWkg1hZ7SKh3XpP3QnGdvx6T+Hpu3+3Vf5TdA+gMzgvGvOtPAZcWXICX0w1eI
cWV/O0R92dmj0IfrBLqOdCU/jtcoV3mF3NZoiWurl7CxGmJotOwj3X5rnT8ZoSle3OJL32LpXehX
5w47RYK4jyNkZS5mrziRr+Ejry9PFkxn53ND2H4qzsIH4MzM24dTPBRolj9PIkBrwhGo2m17t9Ig
GIFo1qBgwxLYr1rIukNa+9zH7v8xMUXFKiqN0PSl83iI06G3FlhLHiAvQXhcKwJgPflp84pdqNMe
U3mhMXPdDO6PTiabCdGXL7VrCd9Ba0urkaQuJ/CnhK64fTuFSPnZvaXxUCCSSjLlWgUESDpZVpk0
fhLQXxearYiWPDZkYRLYX9kPj4nSLzQpcscwZXSDAs9bkPguTyr3Wes6LZmYK8UtRM6F618ktYwR
vSbQfnkdTkn7OntRa8BXkW8UOBU5YD7TL5nbG1Je4RwpjPii7axoFm7eOMsrHJ6FBf1+bUJo84XK
g61f4wOZuxLZPI0fuehb40mAbr/V6Yz/ngedwGLsSS2HuzRqdVw6RZDOWNK2Xih4PiXI7/EvLijF
qrFf2r9GPdp9gcB3O7nA12lRr3WWQRStrjxIH/r87mMAs8aUYNHyWxjUL5Cj25c/llxX4kExjB+s
Xzp+W3lFwHtYCMvhqjmSifJKUGLkSK5Z5UGNerRCk21+6Do0g2Ozp7ptwv44D1vZYfJ3ZQJCvZ7T
MhHLJ8+92u+3EpkxgmxHwDRUjlNOjsFT4nRIDomLwgm5hPww+/FA3ooOwgmXZ/uA43rq5HN4z6W1
U2h8NEUxk62ThAD2cV3NvHs2/6cwUY2cExxAQNJwpl1zWr92SGFS7s2l0B8kO0LfEMajxfQ7N19C
zg47SQVtxYFw5WTeS8ZxDZCAVQqDzOjDa2VoR21Wfy1S5bXUcZmfsiAByJUiGdQNDWGQ1pStg5Qy
PTlLIEtM335Bn7vO+A2FTU7qaHJCluQaySMUGGtQRDNE89DZP7cKj1HsX3WOkv6Sx/O/u83+TA7u
H6Ee0O5UR1F8gdLlJNekC4yLHAQ3yLsU7ymmgQGQ1RfVY2/Qn6Cx/3hHhaPvc9vHj6xfT4k1TKHZ
bdHrz18ShFfZGVHiIsQO0g7uAJjrtKp4LaN5sLS5bbOZLdkvmuDV27LtBqCOr/vhr/veIhVSpQpG
PBY06+wchM76M44VveuWdnIl0EKBPsnvAtdbP3Zz7fTJYNgrvJ6gX+j29OZqt+JkmLI+q7nrEXll
pThJ4RFjjUw6HwpnMoBgvVtjfjFkyvoOMOvU/twpq4fNb+AIss+Yy9IZ1DUNt9moZdQf3UHcKNpU
YyJoDKvazGZI0qPpj62sz4udCepaFUi3fcV3I3OAbq5c5vns+g18JmfAIwdbpv63dMJAhBMrPnAZ
+Xp3cQFcXmpDysbBJTHjAfwCXM3KXiQlfNc0Xp/2SAyXvbKWMrhZ0YPVGt4l7gYiQUSOBIfso6fK
ceDZGbF2x4DwNxyyP7BJSOsglPYDAduPPFNIdqpOCNLxtqIhQ1V9zUYAjKonndplbiKov84X/Avl
sueB5JJeOWDvcIwbnk79/A+iUkL/s9DfBokrHQ/Z0FmIWuasohJSA203GOgI4XKmTuS+JEOkyE6D
l+oDdWoEMYC0nS5B7fMM+J2Bh8/ue8Ol1vtcrMKASWS0gX/byEy9EVonccE5Mh+O4OUTyds7pGQg
2fX40q4yOPEPeOllBz8rp4RoJbYCCNyzDih58D32r+ozfd84Bg7vfMpGGD9SEBAOHZA/pKhZYxIG
Bs0ppr/Lj3fGzgqOYXJFZcQJyEi8XleGGa5Qz/wKnRdSrD1uuMMfOJ4Z+1j52YWAwpETzM7naGmH
Dcmranu0x15cXVi2XNrLcnc3JUyctBwSYrkeR3vLglWzYbdRFMz3GnftN8kPlUSOKnUwIYvE+2ID
pvxr6Ymp72I/9Pn/GL+ReW2rp6zORnCUhSko5liT9xBjbbQEIhJKlrBZDTbMtlbNB0OkXIPwDS/T
EaUsVSag5cxaA9uS29n5LglWjHkp/KsGf+uNOFk+CDsMNlhfOCMBZPgZN7wsUQ2n4kgGcprRQuIP
aPK8ngveAr0p/o4d0Q4OCPBl+e4L0jz+LRzfM1ijDyGFxQc6GMx/SlNRVXiszWG3+pF+rTUxfPhb
ms4gpMpoxOdTsHQb5Ktpxnkn681d5dg1R3ahvxkn/l0CQmjInSXKm5VJfQZEkflLlsE8GHY9lmqS
6FRtc2BFkBiFqQe6hu/U0SYSy1p8QOt0VLj/ReH68p2943Kssn1j+oZ/CU2iT+T8vgLMYXMYz6y3
7I1lBDAJwcxYCfWratp58C0/dxZBIbf8tMW3if5D7RnQg53vbiujLYttP4yktABLU8h0O+wX3zKf
TIMdTZsSllxoqn0a0wcmBUjhNXKmi41lPUhpNFntQcMn7kpXfTcu6AUMuWjRJxG2lLvKULuUPZmU
hb6IwXak17tnuC6L1DCk2V0wa6t9TdP6OcpgRc3/wbAJVHdkcUDlgNSFIjbHnZ79mr21zSfTBPmR
R8/9+vflc+y6cRIprKyQ8AdhF+/EfV0QyUoOmu/VNYRdNi7HiGrSB20sg6KduqEjxRCjZC93ha7a
/89YER1zUqePC/g7Dz3MG37Wp6BanSiLGZ//lrXA+KYCLCI8rQrmpo+upXzRJQ9Dw7V8U1TytpIe
cu1LP+ZRxTc5VaN1EIev2gdSjrqJDb3D63pRrVsPH6/apgDJ48QdyPPTLTHqr1BeC8LYmaD/hPLG
VoolqCanZBW6A7rJddcj0D0xPTYlZ6dNLeqViSt5UAWuGydHM1BpjhYhz3QIuOKhSuBsr2yJ+tVB
Hhxb5Ewg80Mcu7fK+O6j35DXJUmDdsqCZm4z6ZLmb4zIkLTCUInSEmo6eJSH6MNBQPW9idnhpDR/
+NL7m6Ts8mW0JFvhl/dkxHuZotPyaohEL5XkPvC/qj2VAeyaF2zWbV9thfd3Om8G24105mveObhv
iT3hjH1HBXfvjd+wBKtkNvwd8RGC/l9kKFk4JkYABeWWkZ/sGAs8hX4rzXYslWB26aXPusOXXrBg
Nbho84YEKQnN9lqYXiy+lARdPNyt0mcGiwrnFHnR4ZH96abIvla4hAJ5Z5ljdtquNRBzkRWGfzcf
sLRdlsvLAgX9hqVQlsCUL8L0rmjbDDuwVjYVlietMwWcjE7bLD65YD5ujb1TwY2S0h3hNPigdm/2
hrRmnwqC7SoQAxI2/v3cBn/MqMHTSo10C5OKuwE3Qy0qP3C448BzYNS8FrCcDc4tdDc8nEG3kqG/
K6YRmK9+Chr9frgvfx0rP26rx/1d1BOWSUH7qS2E40uqrjP1CzAq0bC0qW6sgrvx3EtJSJFfbJc1
uhtNfvXUBU/iYJo1QymWebLRjBLBZgTQGyGj/1KaiPPADwJFtK8o/64nXiNrlwgHb32Pv1CVslp/
R5xSPjEvV/cBSjBaTCi2NEm9/8FoBoVgi7C/m9OkteawcbV1J8hC9jb2zr0OdvY7zSUPBJaRN08d
uWfsMxFxfL8s8TpoKC57KDmm9LztlgbQ2rbZQDqZi3MEQxAMWh2so5garDwtAtYKQ1Kew2rA9eEh
3Q2/v5O7OZ8hni0Or2+DrK9Ypc71S8acHFZNWW1vdj7C3CRF5PYZHURfOyUES1t2J5AK2fzCDsZS
DmyPx5uTBTFCXYjSFX/X71jIz1G7EUmu4sgMukoITGdBJT/hhxLAcUwZfqLiKsKwSqdPX12ehHXJ
/M8+y7p8DPyecRV9cQUkXVihKhxCGGwIVEBh9Z8D5CVWDe4pkNU4RwYle96fLt286Iv2ungCLB5T
GhLq+MxT+TfBJBasTyZVbnOFw0mUq0ZkY5nRNm261kcmMyACLEMoij9U4VWCvze1/PixAnboFUnx
5obKSIlHaW5wPxwIJu38QNwVWm38zxPrd+2wqOpGYsf9CRxM9ig0IKjbyILH5l9W0/bcjFHjzGjq
SrfMFwOU/+KzqMNE94G1/j6C9JA1UgH3zSKyLWOrBeaT0tDtGvsH720Ywbwp5khRlKIOppujj0K2
UUTjq2bZYT+cGsuJS7VG8c2nx2JhiQuPTXoJqzX5LKXYf5XU8D6ZrcDIeTLE3QLsgIr4HFcltgXg
M9P6cLMkirIFnLrt2JGaMF9s9cIG/skNzTseij0VrdgNhUPCgwVlNc0A38Diy1Fx3sGzFsCVBdx1
xqDzwBhm+t3SGFxOvBv51oa8BvTQMMuRZcYFBcntVnGK7FYgxVl3UPOuRCMq8i25ygTy18av3V63
GE0tf6Mn3jEqQtS3MvGY7uGjhx/9eyLZWQz/Vj35B6e9aQ4a1Mx/oTh/NGibzgtHrnXtvMAaLB4w
6sMkPVehiis8wUchlFD+hGYFxH2fEq91nkjNJEQv96VXVQOHCj6qG037aU1s3pbzIngVKuImDow2
8ckSFw3Okw75a20ieI+yjcS/Du2OyVQ3Zujnq0vcUgRnaOtbPhYwDaAY//lTGVs/weS/GmBX4ZFg
nta04QH3pN8RqiB46dYSEgXwVfoqjvHHKVDrmtwd+J25FZr3uQoIqtuIaE+eG+ralEDJigEMQGl4
elZ7bSi1jF/08HYFDOCg4pDKb7HA8JUeE87vvfcuY0QotA/X8bjFPBy+7VqYdCaZI5J4Vig66kpV
O3uhxwUIsVzRNPGDUBcLGUPKwS+z3vx8EGNlk7PpvmpWK3Rkheweso3hLEJ8bK3hVLWtNL+4tatx
yJUOXJ9Ya+bfSUIZgsA83ZEBpH6aeN58dfC0DjX1nRxWGr1r98WV45uCsuEeu2CdHP493rW0/mLY
IDGQfSntPgm8DE07UhedgB2nS54P2db1Sm+uJI2tHYz+Lc29cwTYfJKMong7RjOvNxXT44ZxyGbr
ZHVAg0SRcu3XNhdXa4nTrx6C14N/5wSnK3HNcekpoZ1VFkNQrdVypZxu9QueMBrDEtqnZkyioIlh
umnM+aOVXz4Rkr8r5v0kHmPvnWGpyEyutjzfd+J9rJkhd7mQOR84D9QDuTV4JmKf0n3X2P7MaHRH
MMdk6S7AtD6qiYOWg8+yrpke637aTEG7xLlG2eXAHf9e9u7kBv0NqELPfBgaFLoVbmQCuMwX6jo0
GM87XeBHdFUQ1Ei+HLeBDEF9F/+XXP9zvADiuAuvqi+VpocsMsESqmt2tGzhXlGTqPv4hNNED0tq
hbbF3qrRPMPJF6CdQGlUf643jJqsgmMD+NaqU1FGQM0NCqWDhO3Vs6tZVe29xK/pz+AXCUHUZcnd
t9P7wW/sJb2H4r34FY9CUxiaWtrPWwVUtdzOQBv2vp/46CjuHgC/l0GapomqpftEn0YpVf9SIrYe
Ekc/XxW7wChro7RDsDNeD+RzLIJSo4+E0Odov25a3EyvEDnGmqSrIuxAARGj5nbNQQJbxsHeq5aZ
GgF8rUJuXXF9jIL+Gx4sdgelG7sBxQ/nwrSPEumzB4bzKBqwIX4VEZMunwVV9VQGYSRllJ/8+D6X
mraybEgLlRtrLZ+w9VNICn4Bn74v9fltCTtlATeZQfocqfhx/VrCcJbTmpTS6d1L0xOY823NZd+r
E9PKDKRt6a6+R9UHe6f7TQiR3oHnwb1IEH4DGsFc3776RmENrriW6WNw3nCAKA+/1PUlhGoumO6k
GfdER2TKNIxVDRy5O3ETl4v5gflm9lLL4yP4TAHAtSVMEWdV9lv8iFR6NQWqn9yDXotYklAIZkdd
1cR7pKVU9wZ6IAX/WbsD7wns4lu2ioXaioWje5Ugl6Rmu7s0If2a/s4By2CsYGvyjMPwH6ISArrw
WU+0ORD5lEEc0B1CxQOjHlBQ1ZT2rtGonR7nzW1Cz3Mqawt6oA2xs87gWX+cEAmqlyONkKqZ2/kv
qr+XRYV2deOFNCOZ3OmO+oLAPBLKtTRZds5q8wA+VQOuwjnHxfQWZDgrYyzR0kg+SZmIoxHkMQQ+
Nk6Y7hvR68WCZtYddH2iRNTbPpwZ98fT05+sPzqkD8DZvq59+kqVHxeBS8w1HxrUSCCYrZ3Tmitt
Ltus++VPG0LEqk4ezHJRpWibCvxaJXvkOi+oU5f0fdiy2rQhZeNPudkiMHopdcRbVm9n5SaJcSnq
0Acy70ArjRANxzwkCrpWL0FFsWu4YZhd/DwNguH6j1eI5iOwvzG93Xx64liJzPafOcMb7xBlgb1b
ri2vlkS82ABsLA6Cj3Ku6Nj6S5KkoVE5GmjT9442MAgDUdjKIbZpANtZfBMvPj40DXe2jGXBLvro
tFHfOi1LKTJxg6CsbQOksnh+uZBo4z7i+5op2Uk/l9nK3AQgeWN2SEnqlIiLqab4zsQG8LtTolSN
n3FivBVvRl5OsaTqn8VWRiMfX/I+A2pKpoIm9aINycVpBlYJtFbt0EJBsDNb+4wdSzhfEDd2kcNC
cAxJtHDg0yrYg2DHTpcHlJss0nm+YaA79P8uIzvhcyuwl9OUlvcsfJ6OSYQTwGkDFANX7zddl5Xo
B+S6f4KsL9e0+/fRNy3Ric7KUNLFiHE3dqu0/CMkl1j5CE2nN0IFvkYhEDXSxk/xOMXY3bGTCQAW
cjcsD7Bsq1ya0bnDBICYuk1kseeqOXhDuedtzO9pzWHBVagUqEHs/E2hHFFgN20kmjhLOtHAJ1KK
QJZNHfKyiogmHMH1dDxv/xbmwmBRc+IXyWs885WH+PEe48bopjphQNz4wkVpW34av75xGT/x1U+k
2AmN17NAGMeRvRnc+njdtaAvvoQnPEDyv5lMQnBnlfeZ++OAoBC0F0BNAtMoxKCs65O8HcvG1PBF
BtjXhD+Vlq1SaPDb5Rquf9epadM8l07uderculemvaGF/NB1opJ+0HMnU92giVnae2zSkjMOA1ar
EThZb9Nte5SpdJ/Zvmjn6DPi8lSnpw34/ALLHx+paLw9+xKMrmViEwrYc3jNwnXdW5KiBiM42Zc0
HfgmJ91Qy2BlpHiPmhHGG9bOOQA3CZDx/DLw3PcK0Q/sSpb+fDcxjVcWCw8TQ4NJPitVeNagmN55
5MLq4OomfX3o3lNxIHGYTN0NaZgKRBSSjIXvp9kblIjufP11JCJBLvKSYhf2ytapVVH+wZxxDB5m
VnkeQ03r6MrA1n74K9uzE6nTKr/JJLS5+z3iF9VqIS+yZ0VWllj/sfNLj22HDpyz/4dstqrW2AOH
aXOlWqydybcrff9vAJ8EfqflbdiNtz7Q33ynye/Ey5a1FlqKuNPeC+H/bUQChbSgqa7RS3PegTgB
WjFI/++uReSUKzGdWBl12OV4ep0GGixY265NcGoNHfcpn6TH7nUfVSGz1yLU1D68YU8nlO9vCUBc
b7jdUOwYt4TcobkBQS6bda45qJXahCMN5cIJC+B94bYx7OkOxuoZypCuLhSkt4lX+GVXdrqQML/g
mU6+u+R07mUeEiPG7YWUkvasGc1SLl/lF5P9j8UlFikeAk7nTysZrjV3U7q7ow9SU+q0B74pC/Ee
4MqUhctwSsnPs6zfuU0pyenNrWat7lO4+XW8wl1jPl1aD8BdYZEhOYozwMOuWuHRkFc72sxp/OvG
7rimF4Q9HYRKhUiUTL5id6LuHlc/G7XgS+PE72H/okQhg7PzYnEzp7bZ4DLJqMa3u3aRuHUG6mPW
OvAcucDJzJROhY/zBfOpXAlNH4ErxhciQ3WmUrTV4Xwnl+vqvb0RpBRzn3NZlKM43KAdsLW9kHn3
8ISGaoO0YEl2jYTsWb7KNcu4T2zv827CL9FFC4KK2G8OKFz43v+QbC9D/vuBtJjTvkYHvEItqwx/
gkUawXCofGe4ylV0FWaZY9iI4Mo1PoA+I/JTtveSx7XZLY+L01XTI5SYACRyAfGEzS7XZgqcXVF/
+ILmVLfmLyUMnKoclVq93qDo9iZ9WCVFuNP8P+d16dwJkFybZQGwsM9T/mD84JQ1b33cDPaOXZgP
0L6XqU3kQ+qw4uZN2U+7A+hW82DPdzmLQifXTNcp4R/ONypPECFCFJkQnJ0vA2myC+76Q96cGvCT
h2IB5KxltB+xuEE/rQJeeBXgdhxJwUoqcWKyPTzqBA8JZGFgxSJKuklgLE0FNAXvKEM0nvodVzDH
ol7joK+G2nMarltyogrwk2UVIVRMPB4Q2y1A5F/maU6N+raqEcG2H+tQF3YsNiGO5qV7xZlrM5Cs
04nDCBSX7foKRvQzxQAvLCwHg8M34q0Rx+sbRIcz5B76xC0uhEkSOryMobEAvYvKWiF3CJinqHjZ
ApkBmxqwQUGoZ3pRSOIl9f6HoK7CbpaLXIqGU2LtYQ8RVIEO6wsd6//n+Y0N5rLz6+18K3EqPHrh
izCtz54QtaK3QW+ZB2cbvze8EUET4ILkPuSx6aW4CRZ9FWabhc0Lz4O1+KuTFlc3pQt1TXWR/0gO
G3TP7qvsa0mP9LnILpW9AWlFVqWiFV/K5BqWUiVOhgqEYXzjrsZ/Y7Tuak7UrIsUxCrw22AyKhrf
NYpWkudOR4j+6xdVt/rqnb4L9d/XpzM5xHC9VYlSvv1jwdYPvj1dkrsWniAR9RRj/f1MRhgIyH5D
nw7K4SffybpoCQB8l+7GjX3vgOVklzj3y8+tRlnZd7CHxhlpquZ7Te7kc1pVvAcqR/s3xkFQFxLc
R+RVo0eTKAzT/QfqjGW+SGkV8EJP4UkK0wVOK0GXwLgC/TxTpQf0Q3g+XOt1SrD+zLkxXlxTUHHB
AWXFRG1/5F1VIPtIiqKgGIyBZlT9O6PwUhCzhfyBd6Xpqf72z+iRz6uJCZgJ/FNzgPIzLnQxCxx1
OX2NQR7G4fMevTMvEoj4ghhrSOtxORi3kgyqSUe7SXv5BvU2djxmhcBPeh8DCPdpFRTcSNpS4c88
XOssURWd0+FJnIqd8zH8P0NtcmHXhx4HoXP9eHpQW7Bq730YPDXPxjL67TYXbMnlcT6FMSjn/k0c
8k0rH3A7Ht5Z4s9v25VbPX7CuVOK3oo9cE65oG3/+q4zuJOxcmBmIjL8DWXnc+HW+PlVaNX6lDDB
v+1PMkQ+FtVOJsG8vo2jHEUboVOgOnaAIFR+ZPMJ+LgExLy42FY2ZWzA+TiTO0e7irN8GrIlBHsX
ycGc9Jvq5ZFOt1URhpmp8se3+13kfudAsJZvJ6OYkNKpKuiXVBPYiZfmIymBnkNY4iFD9P253tyQ
AASXk0y7kxlVYEURiHVf4sT+/mjJbzBzB7gWjzGNQFU3B9hOC6Fmk+LLc338G8ZRV1LDsLZoYQCV
EmXxzAKcbj2v+kI7NFZnUoAAlpiBFoMaGWVp/WUOp+ztJgneJGcGdjOm8hAp9OXdRN+0aea16yh7
mzcP8/xcKGeQBQlNu8b2d/CK9pxiQgNapEjJYKIlt//BzxVf5kRw5irFKh5KXZibIVSlEtopyn7F
AOKuirWGQopDAEinuhWi0vEU2oq1fBCjetpUFBoLP8ZKuvQXcg5nTKgj/PdUWCvoGwNCg39ZrxdW
Ksug/TVTIh1pcD28DuU3w2dfBPldnzg/81/6WNXElhsQ5ttQ/qZrQg79mDsVDnEoqBuGbSpkSYJf
lCip2lICCHNWMsdk92GIYwGU/KxbyjGl4XiIcBJpiWYBYK1whshwBTVRZNOQl7RhzwsQ50ZQhC37
1tk2eeOaz6QSmgsrelNrWOTXih64aUodBKyMbW7DzKkFFHaeprZrhv9dwo+msTql4t/E6OsNgXnd
wU/Yln5bAAL8NHCpenU7NCWktBg9DkRi4X3rumb0oH0mhWIqlSTTNAZq2QsnY/ENVg9gQOe+N2Q7
et9KkGBUCQiXK90iQi/mpm7w/f9Rdcm3p2qlcIMaCnfrgt6jGMB+eSu6VZOU3BhK5SDXpRBEHa56
2AmHcAn5WLeWKgElG+TCIuy7TEwNZO0SgbssSEry/30oofTxLCq2fpK7R1rqnIsbN9Muhabe5g4T
E3whNcRqebyDbfTlN4/FsVHKfixWc136WpoW3+BE8IXG+yNcpHHxHNOCGYwZQlzFtyN6XQ/Jn5S1
rKDhSyW3YTzM+4hROYiVSG0xX09sKx9Mr+lmK2Fz9oOjFJlDowM5x7rmtvrBCPSTxlpwt9RQukN/
oQ8JecW/anUGZSURxTG4eR1lPDfuRUAv1pqGRtPyslnOMZ122f5i1T0jid2XDL7g+uusnFMBxvIE
blKCwM2wAMiWit3tNCMgpH+6zHp+c6uEJssHaRtqJhDiaM06fke9LbASseDNcCR8upoGJCr4Z7sy
QYVwhRLst5w2icOaVoNmHuyE/pWnMD9abN7v37IoB5tdHK+GmlwBiA/1DrTREto2+dp6xo7tNi4H
GpWfHXJypgyjyhoCsOdOArtWYC8O7IQpXr3SiJzKaR9QUFW7y7RaFb9ZGRDs5MiQxcXrX9bDNhrW
bPgAlpQu9kXO0k5ok0PE2+WD5d13YcaeJzvd+J1plRTjxpR9iWrTHh4hvbDiHroUn5ur6BlpFdcH
9yu2tJ8oABx6ZBcenTf9g2xrfNnru+622BfSOJ7JygC9PF/qpAMEd7E8wll+i9RKuEI6w5qyjZHD
anM4gi+typQma8OGkT82SOHRpHq60zXw30ZuaV63rmCOqKqvvZkcTV5ZrSGcLd7j0U/tBR3/R6BN
F6a0QlWOatKpgKVObtphAEu1uwMX9WY37Ksp3wLdHIKNCcZHbE6Dtimp1zQkwSRPMsaVezAfWQG9
O5jJAmT5s7DQ3nmv8irEFPKYaApFZnDSMiQBV565DjS5YIXee4vK8pD/lMknaJfZp/Iq1Q37Ltb1
l0A9HS88+w2qCAkgG+yTwZm6O1f3iJa7R6MPUudwvg0xsUsozuCEMVQMfwie0hhcprwgu9SnCrWm
IETGC6hqdpwTD0l9ijCULQRS9W7woooC3GzsItFVzAIEeMEgLIDYygQfCzh/dd8BWkes/eab1j7L
8j5D1sgSgLVHauVZZnvl2i7nCpqTPAf46aTXt6QaI01jiluQPNmpglZy9NAXpoi+lDOztuWlk73d
1mK3NXzrcqM8K8/u6mcmGE4gRlvYk7bxbPTQ4PmEUHxtKois3dLA4iiYLWDLnLD/GCXE2p1MY5jI
Em8KTHl0QYMUpBm4fBg6XF1lXa6McG/WhYdEjvS9YvpNNx5R/5UbTyk5kcM2vDzJYeOeGtfK/l39
NeOsyqGdAnCABZRhT3TjbQe55lh5qAcS1eQmgbv/rzAtLY5qEDAQm3vS7BpUoXWIwu3wKj9BcBLm
aVt7+Ejb6eVOerTyb/vyr3EctVuRSFpGTtN30XYO7Zq5zg3hW2iSgnb9EAHp7qYvio/IbuDXpd/N
ufKyk7FtA2pT5Cq2/rBgGKBW4WBNEg0sKPxthQzKfFaykiuoppjXClaalCK4NClwkUo5wSi8jStM
hwGhWuXA7zAn6k97YkNr+gln45rNQHYyTH8Fb4vitbPclGgKCX1GSBsMPG2HU2E69Xeq2tUVmO/+
Ll2r4N+w96Y26S9xkXWqQgNeEoxaWPkg1RkIAQemhFbWjcmJSIStlD5Msh42xW1/+iN9uhhdiCaU
kciQ+Kpi3xFz2JeGhhmXhQEKp4k6oWCblN1UhheNdL2BBJOlf/Z074/j8lKSvLlXXXgDn6DJFEyb
/D5tQ4n0Nj5ZCZ30RKlJFHletO08xNdwc/n01NJ/62fq2MnR0WCavHP1YK8OeMJ/2qML+osHRVAu
im/qhTCA54FW+utSkMCWYpbAn9qpICBkPNN3S5M6bSwQYffo8T+9Ymh7j3W1oApVNcewhpAl9kzs
KLMbbP0hzPY9pdsPbPNmIeiD0gnGR/+5DOKOFKW3u6b5nLpfBqXgJfWPyio9yQT5yNhx1bBakApw
99VXohioYVWMVWl7pZDZW6AMuEyATLpMbWEDAnyzt3jvKTlz6iI2AwpT043XSYRzltKnRWqVSDjx
jUYQzn6SWrtN/cdKAfX0fwaOo9twNAkITqlkUAB7Mrzmd9IwMxZYK6SYJqYmDVct86wjkGeyIdF7
h1QUfdzGqOiIaKGhj0onK/zIBT3nmiXNNMNggK7qBVXrE7TrvbAz7dnZfnVqb/qP4lL44syS/049
s4UbRBDkOhB8Y8yUQ3uDNX1Z7MqHS464VAG9vy2LAqgXa5/PkDJ8HpdiSf7Pce9N1iMXxE3j7dzH
F7Z58ApLocE3+ZendAHDdAlDJsemtKnywQYF+RpeDAEh/3iMWOIFIlq7aTOEHxkXJMRz0d5Oc8Xs
w3wS5r9OGe1pQiGBPvXpQKnqoZdA97a2zrye2wpDww5Vo9HBcSyb91pUZbuF0gPeglO417NgJ1aq
n7h6HysnwcxRNrRckDUL6NjtHqRc5a6OlKoHsUXbdiB2o8Gv8DROzRcJZvQIbF+qCTWz/kNxy67H
7sfnkFWiC/lS06KgYgO9qtIMXISTdEN0f3frZTcObI/n69NtZrQnRgQIDr1+fwk8rKNd9v/vlrKQ
vwuyk07NjnAxYVp8b4AkhwJa3ZTKq/6w2kh5KgZZJSHYOtbQp7WcYqk72SZBKBfnaJtaITzqej7/
um3IqmUqtaIA27unf7KdIE50+QY4nV0kg8FzhKB9N87X5vmFEMV2/K88fidQsK6o6DvieML4sSCC
zbnkJnDaEgrNvX/3eLmwxV94UXNaiod3mVJT36sY1gbGq7AbON451aj0YU8bNcosSZoa0tgFcF6u
82dFOYC/zBQSbIgA/xNAN1KDSFBmtt819uFxLirXSFCs0YmEpIPfq9gLYFSvlShAPYN+lnGOhpLa
PTZ9XlwuuVXDJCliDpxD40iJL0l30zi/9/WPnHugVJ4JjZnkNFNPmrkvCxCpFd4EcxudC1pNmVsN
fDv8hG9wnzE13Tpr4N24DwlG+EkygHJ26nQ+5BxtfbsxRBARfNVFJll7RRNm4ndGaIwxVTJ1/Kya
Q7oH0YY724pVOwtuNLjGkO3//OcuQd+YeFBZIV3zTqif9KU2MsxMTN0UCxUtL1o8YH4nhsjsd2Md
om/bIvM76SJtJGQXN+Jx4XaF+rn29S1aP42c8pc7NLjRMY/c6f7mja6DHkeND/8uADAqDnIEEHOR
ZbeoxXA9WQBlTYQQwAcqxmrKbhj/vPBwLq0m+kILCnZFh5OcWLtM7XmKXWWjrRXBW4Bk4eVfFcIC
czuhl9+lMCtvhfWa+6ky0SAy8CVnEYqbeKic4jAoCiZVn2jrPmsAoL/tWHePU4sOsB4yIb6rrHsI
2n9zv+ug4LquyeA4E+Zy5bQhLWdCLawJwZSN/Ac++9T1I4oNVANFk+HddEkzqUeqUdMom6aaPh2Y
ZvAUH7jRHgAQqvV73X9XEL+ZzwkYuiOarhueyKn99L/1DK85moJjUAQLLangAzgXcawaKZD/7kju
UBMoo0HEyixRXji8Ys1Xb6ItxWhjUAuCgEbDWA/7TTNbP65WK+dKdOh3DVD/QgsID6kEqcYSDiF1
W+zImLvGcrION04GKR3ULDALDsjxMpC9TcD4UatKEJWUukh32jrHDcBjRY1GHPtDvTZ0NYRn3O8w
ZMNFXSBcEdAHjO7WpG4hdqYRryH03GCnl2ZzMGa3+ZxP7aCC9I8eTqIQiJizBz/dVrOgIu9vhPv4
h+3nEYuhbMRcEykZ4/merc6YWkgi6lmZsuZQJ9szvQHU2qJgAaiP1a66LafGT1fFbzGurkQdfIrb
+HVqtM8dqNEk8VHBwsXv12vl8DxpTzKKPlcEFCsIyED5nDm3mQonR1yvZj+Cf9XVF3czeOJZ8Nke
8W1AeYy0xS7IxLZsONQ4FaxYBBGWL8JK6KSDsS3UzdV1luuxgStaOEp1SH6IYsVSB8A9q0Z05vmT
5x/sfx9uLoLoExN0YXUP91hfyWt5tC/90NeuvTJff2F8+TpbaXZhJoQq5cYD3bpQbIDthpiulJ5O
8Z8jkAv7zOk2/SEMEyE8oZ8X0eey/UrnwxFpSPaLCb40Wp9aC+b9Q42jGpDeaR30oiQUbmwZLonQ
k4pr/a0PqRzvaezpY7GXXTpUGWGjxbp8JWuyAefbyTwtITmKhfIrQ055m0PEAj4wfYDjT6aixFFr
9a0JSoLxYCzLG0Ols/B32llI1nEqx9ocKKCAFFjOunal4DkHSdAKH7FHIQoTi8BfQ1z9wuxd3NpX
24UMqz4EfU0ay+uss2cHapF3zJ5GKBfFU+ZtPMUE6LjZpKS1cL1DNriVzsF0zxq/9RS3f6ok/n/3
y0ksxSw1B2vn7gHqdK1qAzt1cIxbT3NyrWOf/TdZ5ABuHvi3Q3iJKNph7rt+25wYzAEU03ULggZ4
ZhZHgiKRCDOnm8UvIZD4bZ+STJEaffFP5l2Exw6efnwl6L3484cavI3qM7CjQhuNjCkGPL3M8RJK
xu0KGjFanM4hDJXUL5Rypgapfb7DOk1WkIHSYlpNXfGnW3jYazfzAU3STVISwXhaFfZ5bGG8KGEN
3E5/AmnCuKvlXlGIrews/U0YQd5nfzdf//8sKcAS0qYWJXY8AXpnL0wuIJbBlTcN4aS1zr7bhh/j
fWjWq6bp1chPtSytkejZajJoTbny1ZFhrPG+XOGLRMaCQST5UOsoDIfD7EPgknXBCfkAPksVt5FR
B2zrq6E6WQAmPzJ4ty0cEZ4yh45zsSudIKI5Tmb3scsMyRWC4o35EbarS+D4Uq7dyc9PN2Du+h69
vpYr+24r6GHvsuoBy852DP3/cWSCwFo4AJEAvp7i+AzFzy7tHlQdAF3Kn71J+qw3GEMUiEUcursU
8ZrcrLekWCKDNrb7cJj1ThzTW4wEgtNCasOUeCIFvROm5ENtSPLA9Jo8ctmkn1WS6oZs3zXVKGdi
tDhGjwQUN5uw4Ebe+hXVZ7ZEX2nQxeK/iYIAwtKF8JY0le5zbrS8RDHQShXozRqczsjWUXHgF6v8
G4GBbS0J82FjkbjvpC6aDzhG/yOoBXNdob3lF80BPyJGA7RQxUiJtjx3VjaYQ7W29s3+Y9cfeXPo
dyx9UiwEH7Rj0vlIuMun9U7Z4U2e8ojO4gwwVNXU3MicLsgtFUovXpfYplrCHS9blUDMCmOzI4Tt
IrQg3to2aoPKtIR2wxtMF8d0erOMO2HWAPsuFXaaybM1E8NEbMRBZ7u8jZWZsP40E/3/DkiYyPsz
ugSxNxkYs5Gf98LfFtd4cXcxjcRMG1S+PvDX58mzd5oGg08BQw0Q8a9WYUiwmSGS8fCVhYzz5NAK
47hWzTxE8r9HFMHXT/MIos4Punm4TklxU2dbpPLbnY+EZU+pyWcrBdxnGK0it8udEwh7/3XxdKPO
uI5lNAzsEmysN1DYeOgQ8a5NesqsJggheG9Kc8EXUao9ab5APwxJYRMExipQu0nICAE+E8EdGWak
vjFRhFMR/FSHrio3qfP5nHqzebpHpYOSELK7ZVGIGR4bwF+T2lqb3wZ9kyjCmvJ5NAV73GnGBlK5
kLbMzCxsDioPmPRWO/2PBF4qylVolX/CMIvfHRG7Rx3rPqeYWSWIuPKn4zR1ySlcDjZn6OJiPsX1
20XqvEU/s+KGad3xlpNV4uNqtWnA16AiSlVaBptGvDEzysJ3z4GzAmwE+Gx0B8jfhmy/kZK3LM5E
BnkSaTOwp5AbDH7MuIoq+vjGMXQKSAia0zMNsEae9fEW0CsOMY1vQYrimWxNz3ArwvHlj3Q04cHx
p6k6XFEZ9kAixJ3OkcC5scgpuvTwOdP8GJEASZvr3Srhv3RUKOVlmOVd1fyKUFLXKqJkfA2POVko
WvnsyOJ/+MvlbJjnk8JJ7VADbyB7KmC5cM0ttnt8M7ePFKCIfJD6clyf4DTjl+dwwhCLH0iN2Vf1
RjyWQtIwsMxqfZ/cqY/TAqBK2OJwhv7TbZXLKQpZvwPMsQJZg6D7BDLh3KE46owTT6peMIe3LDAW
LFPCiRYJntAtOaeiWf2NL0ipXJEHZAWCp39jOvgLPudsO53vPwTOT4MLKzSaiaBpk0WOY8uYJapf
HR5meU8avnoBqgftt8g2xnG//QIDYVIwp6OKdIw7sP6wvw13FkcHn/40SsFMacCrAJeeLgafsTzB
RVr+6t9Ww+3Zd5A2CkQwXAJ5sz5b6mXiq+nWSj9vHNRMEIUOs+Zm7h48qnz1VxvG4vdG8o9HUc4r
DCc26C/8QwER2q24gOFQfW4qqgFihMaiO4NGYLF2GutqHgtNgrg+vJ0Am0Cto1HR3seSORSIt1cg
hA1ar2h5vrLugMemxhdyKAgTWQwNyrZmHk5ADwFZiOIGWn7nrO7BNyFPevHeEvbFYDpIBtXWBeJa
BH7hrW4nKSJiGy7/4OFhLGBwfBNnmx1SgfJxi5ccAnPKPPEdsXgIp+Ear869F8XHJqD03oIXJyci
qlQeMqQaHmVYHQ9rz+0uYm3ckbSMRj3evpgvz5ax+GjBVXQHAVS57g2PRAm8/klWlqFDJGfORq/d
kYZvRMTAmAxJ7NYAMtOoVtHmYwu8c04InxnMdcJwNCFivWup4MkZPagcCHJxvFB/tV5s6vquvSvz
rCFFxckkCyZ7gF/WdY0yMlsEyaxmCK01JmUWxGBvtbmDIqaTb7/mM1CGKZo6bZQLQJycyC5EXkjE
JS/Z0rbsqfd+asswYxnLdoM99dqIlsBZ/+/+6TdM7vOk1TBdpuZasK2OdQI6i/5u8GogHGZpiUTv
muB+F70oEYUjyihc1glkb0tPnQdwYD4h+o2/w88wCacp6aNMf6qLg242XB0sF46gSIGv7JIbII4x
pSdblwvyGuIHWINRDKI8zbesHixZCTGaH3OTMdiP4Wld1tldDoiSZ2x3wNbDkCaIOIgNimdruQsq
HGvE25QLbIyHTStamX6tjOa+gV8uUK3WTiZ3znhQ95/xvUoFxGkRh0SreAhydS2P/B7MFJQ6dvOj
WBLUojtFNjI4CT6ll8ShU38t86+3z4UBaVXniuegrNgo8xvqE35n1unrTfij6oHi6FPQ47B6g5Lk
55j4RHe4ktl9N6p9bdB5KzKTOtwAcBTiFzverZf7hhKqqsQmkZrpieROG5bO+hZJbndIzr6nrIs9
vMGbxX1fRQPIB75V0zrcjq3S+FqkKh+fhQd49KvwwgGBhVR4Qu/WK9jPG5tbeTpmCWoMDKu4/lmm
J06J0iPPlIHsrWMbH/O/Mo7Ps/7VnFMGgWN/iMaZn79sURw0de+NpBJJ4dYeH3pKfDdoahZuKMUb
XcH+PjSX0vLEZ94ZVF5yUDFCeujMrz+SHu7+UQ+Mc7u2HJUx2Z0betlXFTKgX7o6c52FmUxggHB+
6CNt/JAlYTyBTBxcvzR6hhN157jq8VCUI+Xg4qFl2lecEY6vhcDs8uQLEsr7e5BaR9hlnV8DpQGa
0WrxZtvz13DdoQ3HT3jo+ZOA5Z4otv1s7IIm7KPtw2D5ffC/DQ7jo7z++gwviVvmM5+zJlJq0IHx
/C6gSaWa/t78e86aDbJWaZth/zykzqd9Zwi/hJEzBE9xXcbTuTgiFLj91XwQQKW9tPCO1eHv0+M2
QpOOx7Hkel+VpQC/BdCDeX6a0rRZZkoqz3fehr+NI2070fmOy1XS6jqjOlEIMLxwvqH8dfaUyy3u
tquGIIao4pl3BCTq3knYXLVdJdhVCSaGiQ5FPPDYnCS+OO0eYxBo0mfEXW7HNBiEpGz1ASA/IwB/
o84srJwyTp95kK65HM0gh21l/vwdWgdYcR6K2A13+DzK9DBXuLXH6abtKnk5FvIdqOdRbPdxMLmc
IHDK3GgUTnbSYvmFqpSgScGVuy7Bq5AZU7YhKxUpp0NfybV+fklrvOXdsHDei2j0i0uyI4JkUX53
LSYiH85XFhpXt8rX0oCNHT3/MKeQ1vJY+P0yoasnuwb5pGxuPjmic4+xXVR4LyvYqE53K2k4i42e
Hj2GGqD8DSrMAXK3erl5gvukP+RxhCGEt2m0XpnEUD1pbSBgArSbFKUzYc+9CLjD+ZQp7GwezamW
5w/fe4ja4SOsy3Ns88ziMmoGeLBZCN2QD7DVEcc+pdiw9kCrjH+S1zW0oOPteg+i6ff/U03XOt4z
4XcMKM10E2RqxZH1+/g1tFXvKevRt8cfjELBrEFC76ZUgQ5ciUyzYuTQs6WoKo14QaAGPUvXsF/V
TufDiQUBbdYQMYKSlL2qWuOhPd5yooua89hsJY9vaDRpFVhgX9udLD4oZtmx1cRMwUbWgzruIHQy
/FiAgFWjmnBfyJKVxwDAf5QJsAi7fsaiEOh9pTamG9/FZTzXCQcJiEcZQkOWKMYgJpoONJ/PxxFR
xzktzYVbeJvI4TmlWaUg+aHNij2mmByif9/cvelu1N/leQI8QQuPx6ptCDhYMIhndjb4aaQC6baZ
bB+EhYche+wEenLmlEfMjIhnqCzyQNLBQE94VOJjCgSXb7mCDY+9+eADYyo8o2vqe5MyWnJ74eZY
cXyd89g/YWcfnQk9LxrMGo/3Kdfv8T7lHY2EUZqIMCKPNYR0961EpYnOpjk0a37Xl6F8kWymnCmL
L1FaUUU5D2Z1UoeOJDPNRGZWa2s7Y+Mrg6i0gv0AKmhf612FGCcB572jy818gNJH1J/6A4IPDrHI
Okp81HdePPlee9YEelwgT02gEfAMugP8S48PcPIUt9tzPpRDT3CGXetuqxRRoHxqccqlmODCeV8o
TRdox6gTNCobqtehbYAZ5agpT1O/gaFP3/oED1DjZi6clc7xdnlq/ISUxeDjbU07ZngJK5eqSl9O
VHEWfVYFeZMXdL/f3ySUDhB0jRx/6x8WC3jWVtWQQn3Hs7UiLNOsT8/kOybrpunW9pIWYA/D2EJ0
SaFpLFJ1UUipP48fl70t+pwTMT92desuxkWI7IOoWWVrOKYyUyUjuCs8CxtxSxCSJjf3hWlf1lOr
utRrT4v2rBiiRtoO/f/xJZ9SgIbfEsicMT05GLcb/PYmjdAaOQPHlvIKTGxug8QaMV7crzQXZvNS
+bHzALxs4xVxyhpaY4H4KkaCe7h8+LpN65HFjT/jntROfqX6FNA6NEzqRcKyNn7OTeY0v/mlNT59
629ohfP/yYzYC+jTenIMHfoDoEomHqFJuGMcYNRnF9IQysV/5uoft2i8y+gPU2wE98IT3j7CVeBz
/ra8BD6SQjkaWcbx/8ru1pT+82RQc5hyvLsVNDVAexWv/JD6yjxYmykAZQf7/+Nkly/GV9ySXyLv
yUZwniyplkMDTXLAZ6FFiMwtSYu9PJmCny0d4SLmijSGjHrECRiB81GtwVyESBZAK0Aepa6Lq+RR
z4kNVvulAJnxZpqw9A05ej+TogeFGXMJhWucR+x/e7vtfdv3zuDB2RxRa5PZXE53uYMcUxP9yOHW
bkVXRdOmRzDlQ6hXyHp3gLNzHlg10ntrOGpFVzNBMjLJdAYRgj4ZKPA5v/1toXjoQQRiM+sZygAD
YXbdhEifYJXXYjr612HTeNnfIZkVuF54JuhunXERqfMdCQkcN9T7iyBxE2mNcZgdKZjfYE2PrZ2N
Va2zb0rhfgLqXgUoB4IYh+ufopfWRG3ANBdqp71UQ1EFP/wH7WL0Y8dcHWxi6vV/Mhvg4IIEbibB
fG/rl4ywu+7ZIUzidPSKcnwh5YPhIWQeQlW+nPPFNs4659mBe31UhqBHNi6Z3yfHWKoVHYUetGe+
DwjMbM4orsNK+Mk6vtWoMSGihAmDbeDLBQkf+B6CKyKNeK1dqfYJQTwnrBodqyB9hnP8lKINKtGu
p5xuAKyV8J+LxDfW+kWEUG5m0FHdiLhXnismmjBq7PMoNp9zEiDeoS0bZ2qlh2hXkISlvoB6tEWM
3dY5FnN+58dOonpJYy578LZNX4r1owoHL+THGQ7li/0CDxk27JWJnhBquNK660bbhlFK7ykkaezY
dP6ou1ouHbxgqiwoe80oAqVt67zoQQo67XR/c0seLY63o/7tTrhesUksEakbXZMYYKQm0ZN+t9sz
F1GX87ANs5e0o7/at//LkLGnrAuHo/mzdC2K5HKscww5Wfo/JCGM2O/nWYUjIDpC2sqoAnBvH6Ya
S4hIDQ2kELqFU3lFLBQ95RAFSkU+100eUmTLeXhIRuWQP/weMCobocxWZvsgEz1jcf4QO+prrgnD
MlGKUN9LZAbr/D2wwC4vWcugXHjgNf/+i3SLYNCVH8EZqCWkJ/cKjl+UKZPt1fT0GWn/OXI989Ce
t9PU6m2i5VrwHMcOjbR7W/7DS4bNl6DvJq9P8O6idq+EfRyGgYkt9pKFIb5ILEI5xD6G9evkumsB
aDdOlZ6XN3vfAQPxDtUoDEuvL7vADIznv51Tr1GGYR9nvgrkuTm4oUU/uKGoZJwE68vHEyDVS9N6
bKrJ8w3eflF88Wey/uAvWhBQ7G++4SjdNFfnSmcfY/9C7K48RK3gJo1D2Rhyk9HDWXo4WeHb3mfJ
u9NllLq5H4y+gyP8QB1D5tLs33tt/VTqWoENfhP8prK+o657QQwWGHWqfAQzyF0EHRbx/emQciRn
lslXxFt9xHNPvZZiS6R6QUAoIWcVcWO1WySEbBgjb3rZJ/qkI/agnlC0q/dKuwk/ccI/CTAPSgph
t7JtfQifkGdfGv3M4NjSGMU7rDBYjuRrlEkbRbdeV7YCYySDk6jKQTqDRzanXA3Aavb4CwqX28A3
AGXJNYeLF6R4SXPKPPiTVKx5lDGB5mdRAdC/z8aN/cfOS8ODBZCnmMsa8EtrPceduJUvV972nBcz
PnBnGPNLM09xXIRO+8aSPfCwOax47plrIaw0Gixo0Wx/7/+Kq1LrZYKkzAlUThymPslwzh5UUf1m
dFABrr/TtWQ4S9kY5iHFrQWGpCkGpYwHQFxEsEMEpJG2DODLXoo/xBScTIGlBGYNL3CXcJEtL+6E
wgy9IfwlNXcwvi2HRbAjmfpzaue16LH4B9a2YukR5CDpiY3HU4Or3ApbsSIYpm/ZfqcBFIoY7vcd
xbr72uheiEFjzOmj3CQfWWlYBZGZ3lF7/7CpRE6x61wK4ewee62nYDEktOikV735Hqy+6g7aPlED
6QrakWy8t7Lv+nP4c5/BaiQ5N73nt9oLV8cH8JnDWzy6kP3upnn0Iqhxpwi8y1FmeL1X7dkz8qfF
WqZf3Wpo4PeYxnZmCrVMW1JYHoW8lDZ7pV7K6LqDvngfz7EVhEaodzsBpBsNavS9bqz3sU0axarF
Yt3vebxS6Il6nfSkODSD32Siw6u3t6jXI4uyhd1jNTfnStCG7msgj7CvLIAb8buza+wJKUcLy0Tc
rJMD5b9SqmD2JxyXTSvuNox9mytOwoj+Q7OO32HJ1wo6uEygrVSTkEcaQ4GqwL6HoqxLBdSWoUoF
an8EBzVHf+H6wVQUUt2pZFgyi7DZSH1Ege5faJoC+KCDeVyj7eg+IICscENSdDmKb1+eYsBMlvGy
AWweUHGEN95CtPx3GDniIYq4Y4bATj5LmLS+GlZlkw4B9LaVeZpowF7c34z/3n3lQcH2z7x8zid6
iHtW4t17JB7C7vy+2T2T18KocgygE6Ds5NFiJa2iP+E7E01I/pnhyPPV3w3BGWwgscKHQUOXcC1S
HDhuU8McWeLXcuTGO9m+ywnwr0K5rTBK+JGQLqJugxjgsFLSQO4gIU1OqKTqK+LrTY1cpdxWC0ZS
A25xp5ugtNtkhmssGAwkiMMfQUrnAGZkhOQ/5ISKvuvPfnvDt2tbeQukFc2U/Dm8geVYzjVaXsgh
kDY3iQnzEczcbsDyc1auSMciDd+WzB1Zuug1yMWL1pYtpR3MVIxX3Adp/s5n/whH8Gnazz5/i+A3
wMtw/zTjRtFf850dT0NC6U6yv9cxB+yWEhrHXrM5ZkNmcNOyp06YY9P7zeR6o75tOmLEOHwCibS1
L0vaxlWQYZphdEQAHHbksHQmAYTh60T9ORgFGth/vRSeAezMAKH7lKSx3CHNMv8g0G2e31XZ/GfL
Qv41uL5BVCbEiadrPYeu7P1sI8/KgSOJwICVN42eFbp4M0tZtWUTukpd9LBtTN+OHONzIgQZbxzV
Txk3szbIJ1Z4/xMj5wS5BSfhyrMxlmfldzrs/6HdgntrOv0jHWuUHRwkpmUZiN9Nqfms9H4KV4gA
i6F7sfiIMJZNk+kjN0DBRBHvNAQ7qLRgFw39QZ3AGZyOp67AFTprLin29dgz+GHWH8zTR+GSqQ6P
vMzRNlWoSPnW6aKSVh75F3gCrLZNASXjA914PaOjkPSAPrneZ2of8hHO9lzU1yALz5tiqAxtNP34
cT14v5YnjlZgD5ROqBqgI0XoCkWF9paIW9EtZzBZ1HvhHkRnp2NW+/LD4jc4aOuKu9Y6fk0hBHA5
KKJBlVaihdtZ7s3bGen1QB9GaxziZ4AgqCobHsEpEr2VVVA09sI8cxITI+m+sGfja1ntAnLJ0w+o
zqPtmkQb3djGnb2uoAicNh8YG6S3KJYK03fgLhhKNG5tiQ/p9T/d94KGnHcE1lGpuiB7CpIyu7l/
hJme5EVRIM0VyHBLLZh6nSV/Dmr7ZnHvXPAmlU8iI0dHznEoJs9e/0ckwW0+uM82ORW6hbsxtD66
YtRI27p13WTvl79rQFBPk4T4yFE5hnMSaspGVvtefOy/FGUIXct4dQ2o4OXowXKk/r7HduhsDClJ
hZcnO2iLvXFy4J/kj6jAgt9B1p+gZ9l/70/1mhUT/tYuCPTHMklseHAGzUKrMlIRB2TOTZ5IQ8t8
6e2TZSuJQl2smJAHrdQxoUPIUWRAOQF1Q8AmqiCenPsYRxr25yZsEcbxccojYrHxgZQ23sP7l9ah
HSDLcUjBkPvbMVmEWzaWY+h02PSZvpNPXtQ5KIQxFdByrmovWVdzUsvggxBYYp65KeCx+6lN6N8e
Q/XHHh688n29SA39LqxCkaIEUh4lUYc1I+1pI/vv3jhsts7XUvr6uWwCDe8obnxcmzpVzPGglfX5
MMNG3urkC5yvnDGEMonFfI4FnMmoNY1ZDfYcYfd+rvGMQcJnP2ZzCjg7WS8XPbQUcQsd4vqWjvfj
/L6ujc6lvir7kYjwpuTybGOL8+kBcFSvfrX0ReqobOlUAUTCBTn63qLh2ei7vXpewaYyhENcxI4G
3syJYl9fuqt4eDOMxcV6A53R9nrPf8VOL3qDyGq48L26Z8qo6QlrKMm1hxfbF75ej2EplJOlcwOG
a+2F8X0XHofZ8CUdqywwCJFx3T2yS/VzEdHV1C37l5Vl67aweF+lB0scAqePIm6PouqMuTgXZFT4
0pZOy2C8AwMODnYwRfy/KA5xG5/OZ60kXWLOWS8Go4vELx6u4UoILEVizAKU506/pDNyWsV+1x7H
+pTsCAJnqIu9CpV1wcI1W03en5MUrn7OW8beM690JX8VfJOsqQGaE/SAmWJfwzRC+22/lRydcLCn
WF7TVkmBuhu2OR27RYeq3ys4x2QJkzd2Df3sdMKfg7gTIB1IuK5iupW+6+bW3Kwnk2eoaVQeRmLm
RgJDpazsrnmBIYt7l6e2g92Rdb8x+QaHk2WQBvuXxofy61zFhtgfbAJhCJNwJ+7iIHZiw32QQdhl
/YBisK9Euls8abdMp7vUNss3+LPLXB6NVLzy9EatUEG+TLyyj+02NpGwYf30dJhSJF5r2lv2msU4
kutdbxkwny7Tu3wWzuK8t8df66O/QDkUDnM/1cBjxGTymDMzSJX0qXAEkV2uRJJQGadd0JZcw7hs
3wTr2quu5mUn9Q8jh7hr93J7c/jx94pTwvOYA7NGC7gJgcbrTAtwixZSQJFzjwMibRxUrl//6Vw2
bLNlHQLVxTF/kZG/Yglmn2EVD1N8SQpf6QCgw0nY44YmgJbQ74ZbBb9VNXvRBdztNesizDCY7yA0
f/2vmKbQICcvtFsf38Z/NKf1H4Gwtcfqelqo75CYDGxMa833sKDLzB/8kPteSWxqE9abolM3JG5e
IJRQUK+2dTqmacJApOn/yXF2Nn6G+qtgLQtrgRwOJrj2uK1OywjcMuZpmOZtSp9o/zBGKgVWWA28
tr+596dFp7i2MsexgDRMSZGvPuad03Lt1OCmDKfBPvY2S9cQbGkj7mrwgDk4SKREn60mpkHfUYaL
UK5RRM1UHbyGF62m3hZZaAjgnaAlMXSnHAr44I714jx1YyfC/2FgV1XMsgYWdBHP7hIEJKKUXTtV
Xcm8aDZfugTK2a7/2Fn5kbZahMK3Y43HZJfRqAoJ/rfR4kZcolda2vNezkb/UNArUyfvaiaEBtnF
giGMSV5H/Y4kM8gNx8LQJMj1UUknEVIXsBAqv2NnqYwvV3HzfjhdkVmFY/asO98BxhZgcagjYckO
Lq/b06nR/IY2cdbI/AW3zXTPBV3ojChZBRh+vL7l5bpECuYihDzwLXiG1eudXTcOD30lRRXpml09
jef//UsuWGdwZ7uo1ObaNWR2fvpCL0Xvl1/JQPfVMb9PbMiCm4+FAQT3zAYy1c2iDTUYDd7EMC+C
Z/3nekhXRh88syWeK1Y5OMc41r0rt+WNvjOSt9tPI60+h5Z8ZpEbarbkM2Aba3Z/giwfQ35IEY7Y
UeQw15XBhNR3pd66jFhs20b5wgYG7343XZxSuK7+Ahfz5t9RUfBHD5fG2lW/0ffhydIp7ADdJE6/
Dj4F2GfX39mC37Mu9HQJgkYoJYYyw4zYbgJRIvY6goJ5tYs3/BA46vlSBGdQ7Z+uUV7EDmUUIFNI
b17lniPJNmD+3hcOY8Fa9uFodZehiUuthtrneK5UZkF4GJAX1JgPbJY1O4q2mjYsKH+BwTLW8CJw
qNtfP5V0pLVvteKms0Gr+YCHkYKOQjPUgWMk6XCcJv7vQCKRkZALWCyP4JPdWuHgJjfqad8lPv8W
t5NkIsmsFaCY9f6ywrEPOUvZAsLdJtaJ+Oj+jCHYmlz8UzMw9zQfzmjvLNmN8LVGhGT6yWY7mrG0
zFysHaOhPvu4c/UVewfXz8/J8CgW1CwhhAxB0WtC2Suf5oA1rOsGLy8wJXgOPL9r6i2TN0c0qXAQ
bWR8YkKIdo0uKkBef7XgcAkcbh1dM23xF1vZnfYpDiMBucS5sVeHhnpR+9HwpDpMf65oKIs26rJ+
nDS4UHiIHBMJQH+yv89iRxW1LzxegAoXBT+8TijXARPkanHPwLHNRc7PBg2mctQuWbEQkNBtCVv0
2eAkv7++n6WMDyiF5W6YELMasmt/cLGz4jJ0VSFIVSrYWy9WiHXC7hj8BKHdcCSXHLGYnxgd8dw9
UFVAIPTDese1iZSLOf6Q+uMCTymaQMEP4ncq6VEC6iAFKiYzNjlcZm87YvxUB4gj2rJuku07FOqg
5tAvk8CE7wHLuSs3q/wDNT89c7u/mmdXescGgjuiBt/2d/YX5SPCFVQS9gy8qYrsM580eD3cySoC
HURnpElg09a+cR5EI5CvxOJWBfWlAmZ4BTr3vWIjeV5hVHY9wrBcJ+kz9JDC/7v3Z4gh4Dv1+XhM
ZrpQk7tYyvuW4kJdZvkPDZNoUyaibKsOBTebIzGvooGuulhLFK+rKTosWdEE5iuUFpECQdjNgXMN
3bsqUxwyu4P/hKpfjGm6yuTZIxCsFUJ5uH7T2IbcXiIJUihAQ+m8V5+uCTosG7dEAAYONu1s4KH0
1wBOQOPdZlcalIhsGVNYqTArdR6iBL45nw8hmwt+hZCk/csHSUqQyfuz6tpJ6LkfDW/l9M7vIkxO
qg6rRBq3po7nnVz21hBkKZhI8+B2gTvjcPVjs60hjMoYVrboIBUqMTDR+r34lY4iOHTrHuNsOB83
UWt6yRpPwSZXMuwW3nw7R4uP6spRSkrg0F79MR84+b3iDU/s7zrmpDmgve/E5rpAg5aPA/mRr5R9
zff5PjWDVnthnLd0zeuJBEX1Rr8VhWhRqwgJyIHd3JnvmAkAZAyxwizIuw8VNSbv8s6GYkfVJ1zZ
OVxe+Sw5bEOesT9V8PskW3ZCZFrw8hlaIujYym16vh61QfxnWrgL1N6TuMBmqlrP4hv0fRByIY6k
z9rvxVind/TQ3NRxqU7caAOQ/jGsER1LcF3/pizN4aGtBslN3T4UsKEF6N8mmxH3iIMdLFY//0dW
skzxXVnrryikzw5kl4UGKYeaGUGvthrX7XVHXLZRvJTeIH+5mzULAIhM5ZLwDgcD1TgNMr521T1p
eMDdLWx8jRpMjYH57t4MQcKGXcz0yEk50CKyeHtDveoSZP24M+Bn/OHDGh4leo43pRQedVxrSAxG
/TfUIwgqJpMfw1aQ2NYvyyoc6QvM3ZOJ4XRz1qDnmj/3WqxCrzM7EjHMo9IB21VHaGvFyPM4b3O6
eK1S12dbJJkqRhNGkunYvHEdfUNJFJxPC+NHoApvteM5S7zGS/KodqLQWqnmKa6Odd9LUe3O42Hr
S/5KNlhOxtkxJSVEpsDoTUWzR4+Wy2J+uetwjLrRwwzi1zUX8ZX2isM4HqVJSj3lSInLDVbS+UAE
U76oe7Ptag0YwLgEN3fEU42l+htjy4CDncIvSQp3utL8z8+y563P1bTz5tHs1BSVyWAdNgsmabcP
BBGmctmyIpogzio2WdCkTNZv8DYKzedurD6JYyFRwy0EVwaUX3oN6+rNVFLfKcof2pCKx4TlKHt1
kq/a91ghtz3oG9nla7WoLbLHsE3OGJdKTcXkB1OGAdfdweruUtargV389dWE3+VPTWxmWwPKie8K
XTqCcbOXglz5SfWHcqi8afJX7eeNLJKCKYyTOAxm1MfCokU4m0d8i5MuB53dwRuZNP7DdcxSsB/X
K4kKz2oG9fJOOpIBLUOqmWKIrGDyAV+8HRwfPs7zmgVYQ7HXW/zEZuKiWXFEvu/fdPUPmNLWpBk/
0fNrgMS1kFz+hifCuDF90bY+b/HlntUHm6GK4cMCdXjdCewP9VYXSnYIzukYY6cEI/lBbi2uiSsw
z+HgeXrwE5P2SjryM2kDW3PmsAxR6gkpRxvFHm8jhLPMQ1VgWppgfm58k7xBCvim/ew69rYpv9zV
eaeXlO/RBvIL02vcK4nVXk1zxZTtKtvIo+Hs+bfmIOuwUnS/prnSNe78/29xV0QrghDNjpSw3RNk
aZKJ7eurZtKZcQAQjKaMK+FfsqFJjZCxbL9SvUu3V5dU32hURPbvswwLKDyaS0Vnc5yWg8oDSJJ0
//vZAemKVyGsVGNMo+cG3wNoTR0InLpzf6MhK/Gf8UnQxMoEBgzc7/8fXBcKZZ/br2Pgs6bH6Ngw
n+47tCN9H8qstwT3JzSmYBQq/o7jYAstEB/FUyEoc4AHoSNNCkg+xTwTCSKi6xADRna6kRIdv5M0
8+e6TtU92XHWBLQLnSqXHJk3S5r1RigBQxcIMlb0f+aJvCW5cjDT5toubVcFCZWP1/AlPQXhukPo
I3pou+VTCdIoJ7ORQYWqgu2dp00gr4QlhufhlbIA8hYHetgqwsJ3IMArtbbt64XRegriV2uMCfo0
5ath+gaghT5nflQhhe3RFyIyQh5XeyywB2Qf/AqI8NdtGTOhPgEhoujxnhTLYWr/caK4V9OGQYMm
+wglS9U53QHCv44GcKcF9Mq6j9txreY5WfBj44mxU5BiApyIgmI18SzeKu1AndfPSYTUuwEAh2FJ
rm/l/TleEfESKDBu/Pr4Y1eSPrAoEk5y3kGiYymdPD5tBGcjEkuL7t847s+QQJqV7gZsOLO5VTWb
7STp3R9+L3e455DYOMXWmYBaooZcUYh1Y+491FxTzxVPAmPLh2Cu9qSpWAioVJ/RjIK3GLNhcvC0
u2nSEiRYb229ADchgSLkq04vIfy9AThp0zAb+ldOftqoSfRagmkO9SdiJi5g/Rdg6VUSVKEsUnXS
JlVdH3RQxHkzOV+W/3ycD5JzU4g1pTLdz9/GKoGzKlvizfALVhSDyAFRnuqcEq86pSezcNaHWcXF
2uTOpS42/8sONwJkUes/UAFgbxaEYVcYLtrQ8GddGm5wezP+D5KfkiI/bq6mAKEeA8un5CfuIoEs
3HNAzQuSfznsXYzuhU+C09b2ERs43RGOb9pSL8082yBae2zajU6WAXW92h69GEIHc9n5F42FrTwG
OvvirvYsMTE2bgAonF+7HIX86unkgNtCY6KE5tbwizeh3wDIw7k/YIZPRME9vO/VWXBcK9cDQXcl
jBsEakPPQul2yNbIkLf061W53a22Pk6n2Oy0oODCs/nh0AvxHBRow8owL4kpgnBjWNpvakC8hEB1
TXC8+/wspmHlq1y1Kd1OoTE+VzRBzszA/rGIKC3PKb3W4O3TjndG0G3iDOU53ZfL+7/9Oud/IWjw
PGzXKPCIKqlWPHWMdzmzHXdHpH6fALp2slTE0mvErPRxIoptBhFwsl+ndUFey9c0ONoALCLT26ji
TUMVrclNX2erakamsmjffRPfQU5EbBPLbFGTqTY3b921QwWTmtDVEynNZsMFTsc92LBIyvor/WTt
q1ocjKZuvb6Hf9c6zzexwB5IrdFpXUkapQqr1n0LVOSYxzmPFpU7L6eXuihKE7zgHXDb6p0JTk/F
oHIxP9atokAO/jzacKeLkjCz8pm1a4oMhPzwGQWBn2atTuodfW7RxGCFSf3Bu0W7SfagCpik1yf9
w2bNot3TeN/WM4azwCNv+nMP/S0JVzgETb1lpXZj+kGSgux6pDnZjuO6uk23ed5c4bVCAacl5PjG
ny5z9kiSL+3sBNrlL7Jt745jUCs2SOCiqrDuuoxMNQ9psWV/xaoNxn3qQtdlWyabH16GgOSVkVn7
prCaqur4xORPPfYjjVvR6HrTAOuGkSRHg/XPIhfl/UM8TV6kjmL/gqfw0sWr3sQNDxVUUbMsaCej
wo2lKD5IIa3gnDN3lvnzBtrDDsB34+EGGF5tiTA+bNkSUVJQQ9UnchBXod5m7ZzMm/FBTIqNMKu4
HXZ+ymUQejHZFYddqmUrpBIEmvvgw9iT+vx9PtAvPekoWLuPKiDrYpia1ZLazoMWLMY196TksPpl
jyLqWo4XdudyNab3oWBy2yWdNb8XYx4Ckb0MVs59wLvbzhYCHY4/Srdu9Q2mmE8CVitKf41HmxNu
8lnNgz/pBaq6G681PPwBHVQmTn23GcquqZevpaKW/a8fQJ7jJXarr6YiTAg41BuktMX+UipX1iHa
ARoX1fHhaomEu4QgNa92m3T/uKrH2yYlYTdfc6WRT1DJ0p3oERTBmtNMdBBGcOnm0qi+1mVJqtrl
45/tuLWj9S3WzW9em3KiIIqr5uIJKukXquXfYm/psUZjBv8MEBIEkP6io2LmgJ93JwpRiROynpFd
/mGpB0KNi3ZAzcV+i1LZ3Z4xwczIGpoh4bHIodQN0OY32LZ1dEXdAvj0iK0SAUtKS8Ou0b8drYp2
dFob2V3hStiwcR4/VA07bo18kkW0rskbx3c4wqJBTzIrFyWAz1itz2xq7kwTf0TLFfQETDHJ9/F7
iEOK3HzeU4wCWif7UoyTIbTqwG7X+sZvTm/p5ow7S8tLgEvjLaYQWFnGqs+x51NHfHLiRAAe9Z0S
tpzv1RD2+la2tShMnBJLmJC/EELWYin6GoutcRGP3q0T0F2/m63AZwgNcbPzS5y6TLeFKGCkP7M9
e4UiN0hlqB6wOnWbf3R6A8dxwyqQkq5PvYRBz94PfzrktdhTTKISXyo8cPwRYUaDYBQDuc4J9i0v
DDcBhOu2WEIwRZUMYuB7P5JYai99x3Vmr3n/Tb4zvbHJ194M8YGX072HIvhuELXpBHtPppyFKFvd
VYia0Zb+W+jR445tBJ0hZl6Z/+ZmzovKjQTYbqsGE9QRV3dHjES8/078TnTwpRyfa+PKxRFv8NmF
EDF3b5Af1TeVOzqOmqPRK6HOr6E4+GK+bcsCOwKaNOw6cN46gHMP0HFaasy1eqf50dRTxAtBqaWo
9We4F9d90XPby0N6WFKlknf7IQuPHtKZaLiCPbB4z8ugy48wnl95Qw+hJsiLPvvkC3cxwAgm1M5X
1a42e9m5XkPidLB0xoutgBKWfK/D1+NPh4MAwS2aMvD30kb8jys8hJDo3XiWHuFw8kKV9QEuG7Al
TA5j2SxFR+ADplzwu+/ExXhXIX327nizU8WIG5DaU0ah+UI4O1BxB9jnU/q/hmFA10ubv1HiClYh
E2VLvqb+6E9Wi6okek9Mys/tZlhg99mM8IZ5GV46Bxn96Zek/jzHfKrxXQKiwHhXZDrybgvfseou
o+uf2RwQHrWXvfz3V9ruwg2a5gtcCVx5rt1cQ2GhPWQXTKYYsKLxNTqUd+EniI2bTgmlzSWxLv4b
Y+5qbgrq0NxzZdA023gG5y2lanfpP1EHt0L2O6lmky6vejI37OiT8mcECNaOInIXgzfIcN4LVMOK
5dovSiLqyivQuSOtMyPdzGbr47o+ULLe+HdL3APyMkXFunq0uH9US/jDjGfKN8JVmvMrwyUmngxu
GD813xMiN+7oMlr0j9hRdO0HPeopMLKMpepJCxOfsg8M2lNWnh776Q/O7+Lpb+PWWqcowy4XbBYo
F9QqSBTmPMwDAWhCijB5VNSbXxSdF4G+GFje6yFIP2Tlq8X68OgytP+n2sHXBAIvwLMCrloqqvkk
TNH2U4AKY6xwkrZFclGKDtEOSUzBggVuClm3L5ItDQKIauJT5Ckmh3ha72UD2NVhs2XPCXoBAGWu
dTTEEk6YvQYeurVKAJrDqLhl+J3hFRaxghWmAfQUNNqvwHtN1CgUD7/L0B4o0iRKui5MkFnmcUFJ
cRJGrRTmvwMkklwmANnpCLT1WZwEiqNnhpXcGhQSqT0FImoio3Fb5T+lMyfRszL+HWc4qUplurSN
4nvfEbFuUEYbeJVShODmWCW9gealOgnryr9vIjnlc9u0r3U744XY1fd6YQNmN2eIGkgTNL2jIc/o
TmPL2+3zFoiV4q3OBzeqbS3FhtNfRxTluNsUYpok2G+4LXT4R/+PWeuVySYnnffpq7eAyWIva5zx
X4J/isHAXm9xlsvVPcIoMlE0l0g5+wFyrq1CV8FMycgQ4WcFZcJ+RNuHv32DWLSTrxKnZjcIwvhL
G6z7TPWjOUhRfAHBCEZOGrEk1B/HRUoCto5tiPXVX/QYHhTliD6hE9pM/yj5b1YFRyRMmFnXMSp0
QGPO3BIFMOQTaBv4rw3H5IJaAlE2sVLKAFoUNgbWc+wbFHrI0BKGeu8vyRg610aOyx4G6GtLUCSh
aB4cwsHtYBPb+k+rfKNSd+LdjOZIjN0gM8X4qWOa2IYCdHBzV/NdSWYZS/6tRa5Rc6XhmTZYpcX3
TVfiJB2tuhSRxjtD4ApmmCvTvMklpMhlI+XzSHqUMKoei2u6GVcSy3NFWnIUWcA34xXEeu5oIZUW
2fWDMsLvbbjRWV3O5j/XO0VEORAFQqu5pnoBdx+K8qtyE4OCvg8A5zC47eWU1OGAStwQrvwSIsJF
JwhPMrquGe+1ASImmBK3OQ60lfkoCEcORo9kMi6MMplHBJtE0yTNwyMKHghrEds5dJpOMeJUt4fB
k7ecP9UM3t0zKZ/3Z+/wz/mtrHGYs8Y3zpTkxgi/yFHoFnPsF1tE/RDqb2UWMxqNbLETLqngV1RE
nLi9kGsJGR62Yqs0kbVoMIGxNu2uwvnvuioYZoB2RAuOKqQq3aHWomdAPA79uUaY9CKVvYPpIq7T
vz9c1Bf3yYrNFDlu1oEELrgyRtotYVSXxHOELRLl76ldow8meMl6KVeNf+DZ5iCHsQkLeDJYRbBU
TJhbwbRDlln9QoTOvlqvCdZDqF40lvt843tye+8iw13z1h+ERvDj6tQLYrhc0xirXNagnmkT5KXG
ZKVc22xvCozh27/1TxHu/GyUzB4twVjDJpeQRTusSB1WP7EyZSIKxb0frncxGGThvZKZSq94/tNy
IIrV5lno9gAS8xa1IJ5XuXISWeuXLZujJCUlxKY0dzMkW1/jjU83i8muBagzhbFpVqzWHE6OoJ9E
7G0PbrVLwnZZeCTt2fiXkQecONNohH9LUGhNyGEAkSXgKiY2RFQWVlhDFhV3R8vn1gDguE2emd9o
ugj0Mgw0QqWPdK4KXYANGi4oXV0mnfQQWlqOLsy5HE03Uv8jGz0rl+0ZB3i3eajIlkjb9Cs1dfVq
lsLNcRdQ9VIlMr45bRw0WGcfqH77s1qIA8NoD2nRkPtWmbP9BdsSPakPnkv46cRXRj/ufB7PEYtd
PNoiSFXcfOjfRTk1GlgnGjwdx59hMg+soVZwetzQTXY/AEv9oX+dZ8N/wcM1tL4yUW8F653U1/5x
yuSo/UrSy25sehgKGou3mZpPl+SBknwCtYb6cw98/XPUpg/3unbXBHMutyVL67EZFqUojSnh00QO
l8MPJRb2SQToE8KckQ8LfNgx40oLZE7IjFCZNTB7F/v5SxZiTEhq3L+Dhtf4hwhx5upxb11mj9QA
VlM29uYjxkGZxgVns8RARYVirV+0CCzQ8whVxb6hwgfdkTGEigT+00ct8vqFM8008Rgd8yPd/PNv
R+rwqs4WvRGP1xQ0YwXib6EliiM4NQgMB4haBzu/l/Tmssusb44wYVqQ+LuIA2cSSVnmprl3HQQF
5u4rx8A3uZFFNLCwsfe5N+0cfpkpVzU9MhnJwCNqIKyRWgPKVoMgne0Mr37ZqcFTeSnW6AZXjfmV
33rVwzzg8R0idj5D6KeZ8nYoyyKdafl2YMjGtECDXb/9Chp4FOtdHJ1n2EqGwEqq3NywnNzx8KAL
QZVd3SMHegScgZWcI6MZmHDWkEB3ipE12Rif0M+yaf2nziECuYkwmW2u0rCAV3oBRLc5zINAD38V
qgAj5NwUDU/QQUWv82n95SqikUjs7kTHFJniq3dDKTbGh3NGypgnGKJDo5mT1V8zuZEKuK1F2RPn
rGJBzNxFvHai0RlQJ20cfjGwmQkWZ9hkMOB0V0eBk9PcIpsCuKvqshHCLFYFEQWNgYMrkZL4/nsC
TbyjOi/z73Ox7CElxgvhvZGxtBr0vFNGV0Bl8djhDL+otuZpVuhEQ1pCo1i+FXUKSl6My1NkWevQ
5uvL4DRwdUPPd7K1EGbn6opp+RrxwoQ9QZxG7+9ZgEXuXHswe/ZFJom2jv0WBssgwSdx42Uri4xY
GvCGio9+7m7bcj9Yxp2cAXCNtCdtJ8f5GfyigDycDPif49Y+xuy56RXt5J3CfqW5iZlHUyCKQQIq
C07GXrX7qsGQW7biNhTiqXsWLw1tzU1XYP3eR1U0NGNOlHjMmUqaWVp3J5i5bcA2hVZEHZqJVpTm
/LrSSWhO/prup89+SmfC1NQ3sdqRfvEoU5XoBtnPSVyIWxXAeWMvNl++dYaeQtHN5vghzRY0E7CL
m20FlelNKLJRGKsXqdXs4z49tSCCniOyZG7C4D6F5K+iSQ3xSRw44yMCx7LxNJNVIxf/jKMKx+br
sZ/Dc5K7ZM3fkDheIAd6L4jgXrrMzoXwEGOf7DybUkPULnsI/TRvKz0qAOaiVUOncKXtQ5zOyQ79
awyGCOjdjLOkEvZrOy4JcvULOcJGQixSNicRVTjEFR1BVKM2WM9vWFTSclfquOZaDeTf8i3mNm2Z
4dwhV8N0fo5WaPSrqgLTs4zo23GreVME7XatJeM4dIDbiRkEn8QbcrvUSwipbVTsbsYpMr43Jh3Z
9kda2SAl+btPg0dW0l4qccx1n8lRFd9TBFNDWWROu2QYuUveSAep6FQvGBSxUuE7EoWmwsCISkX2
pW0dFaXMUlS2qDWHbNWUJyd7hyW1sGw5HYoGu50fFpnR0als51RjK6DDbli6scuCHc8JsHkef3CD
ZliRfz8Kc+r7lLmLa2+zY8HvCKl0yfBztq716Od8vHT2w5UnK6MXc3COCJbgiRWcboMqUxN+hGb4
0XvAlnKpR/Mz5RDwlAAWfWL8jovt+Z+ObEwp4nNYSkv4Q3rjtGnGEfGvuFVsdooG1gOG0kJGsj0Q
fyjtX3vUb3gUa9QW7s0ixuBo1Vd2y+behDASekvZSLlQvABHTXtlbwwfCp/oSPmy3KfU6b4d/cZS
DOb9b5sDoT2ztDD/uuw+osuxwrp0SBKoktI3OyY/vLFm/zehX/KQGNiD0IzFLGHbD5qB4+RmpWuv
E02+kacCqzm8XnDrVn5doUekAw02R1ZKSp9KQQe6G0CULXpSrZSe5rg9+elp7j2zGdPZXtROvi9I
FeVbybs5jefDTr6jW9euPZp8QI5OgRbe4T/dSdDv9MssNDY96ZZGwtMxplkkLpDUN0Ut4kTjxHV0
qUf848awxGHb1bMoH7GoVNXaNuBNT8DdkggI/QVzld1esr88ddDxr20MLQvqwN5ZX+hRBAlSvCtV
6CJwqtWRxPaVZGOaH+RijAgVqbYvrJ8rI6D+p94kdUPst/RybSETddD2MqiIoYSTRDDuYhX3m3o6
iEdRPvlwMQugCo77961neHC2c2xkUy02eh8O5bR0ZdD2UtbqeSflDRQObXwcevxokW3Cork5JAux
vrsL1c6DA8aBIazMweMpHgBGvESAwd1ljdQUHAY+DAYuzQkDAwFyC5BBr86JtYUoN0JtO3wzFCc2
mHc/Ea1/qmYQs8dvgU9qgNREddW/1bed8BOkcBYgZu5ka5Zum7Gk00sFDE9JJAJiUZXJAzFILYC/
ZF5Ul1G4EyShFArSr34VGz65r0vI/08n0vM49FXRpjtLBcWVU4wCv3n4yRgkJIrRDeUbAW1AutnO
8fMsJuTe3mMXz2Unkcnqdrqb2j0lOiS83JmHn070rCvY1oHCFrBWNx58mIGiLaHGLbskYWdLO9w2
XSc7AxxUFBGw5tfPx7H7lns3ylq50l4jgP1mpEiWUQ1nPbPd9gqm+D58goYweHyZbu/nIdRemTGf
eStAPSKQq66dN9M12bNYGKc1ZGNWXeVbUJDLTLMH5Hx0bCjD5yAH0i7UWtEJO4LZNxTbCApj62yQ
xLA3ODWI+2zvXuoAj7rBn/JCRoW7Fra0Z6u4ySZAqafWKR/VW44ymBa2syjrHKhhCAbFZBimXgOz
6KHkP5nvkzxVQZSJJswxTWQp2zpOsVWPNvZ8ItWRCpLzbIRNphO5UA4EX6ijiYCAqF9o/SY5IJi1
5VEjeO2Xa/E8rigfYf0dcLn37f3+jAiT+OSpQOllWOjLTNBZduwExewT1dd26zJNZApjxsVYJDjp
hSRlnSVmC26kkOgxw1+JtVycAHgeYqfCbmfRFQY5Vfa4QEipxsRCZUM0dakN7Q8XBCiapB4xgOH4
NkRuWwNV0TDB+DV4oP8fdQTozWC788+7hMrMf/BZUFg3is5komp3vUl23WA9v0WEzvfxsrG1qU89
x2bRF7vFDbxeWCLGEUI/1JKpb+4Dy6i8nOjHtzxl+8iFW3o1JNdMMWC73UmBQh6af32og7w9wGm0
kFOjldwxbiFiz2zlsYORpqgHgU9PNXEdEOZPpScwQjX14pF4JFwXyGaCkQTuklzzLrhLo8flJCcx
uuaDh4oMWVaMu3fs9jMGWN0WvJQ7DcumAYPvbEEu2pBzEFR3dNJ1WiJ6SBhF/+HmsLgiuUxuWzPS
gh9KAQ7MToLpNcxsPEAeiB/QVElRC1ICCniPY2clbxLOqHxOleodH3GHLom1Bb8WqU1sm/e8IwE4
NCOr8UV8nmWrgaH5o0luXEPPuNAz8/TjtLp6FzDLiZL6wkDluhlWB+RGF7wO6v/mjqjN3uSiUuUL
psNqwCGqcX5RMgRfXZ5DAJb/YwtSzk/qtyXJYPOa19wu0i5NKaB3pTLmbedW0tc4e2DBR7NykDnF
0HaSHg2NhBPFWMZ37QNu3nO96SGgaTDnvHYakcw5xmtERtFAkS9ef27HySNTQ8BVG3J5AMIYCvgx
zMnYDcWS1KjO9JxpA70GnDhAx13eMryeF/6rtWySNZ2q7PtO4MUt5Wwj1WTaYp/9eZIc0NencxNl
tzpPhA8Y/qik+QU4iAamhIJPvG2BZK5Wng4QSZrXGk7XxXcLeEndZY9Ix26A5O42/1FplfFDw26y
bCZ+L3oPTfYclmuMd4UAr/tjdulL895t582CMa7jXiLSJ96gJX2ewW4KHHjvmLYTof21iBMYYQpy
PLWy7YAH+sRN2Yjiif2oOK7koBwj/SFnWLZK+muDYI+jATyjzqYW0PQdNJFZdDTNbvJ1ZC6HEM6+
3G8R82C07EMsXfddGC+LdR48/ZfBt8keh/jcFi+37E1HHtLp3eoMRZcK3IALL+EUkeZ0HPcLUs85
cyfbJdtlEFqWgVhpvrVH/c97XtmXJ7wOKkFR4jC1v5YyuykkEBd/Pu58kdfsQvWhp9N9rRCkruFR
4LFvEtKAX5UaH+gafw0lqyg8MZu/qysKIzwMJKxbmYzpsfgiWt0TOjIph42JEX0IwdWVRkncdACl
BcCIH9ysbW0fPtnhFxi5tBIndsn2m9n4Ph3z6c0+he/Ui0yJirXyWEMZsm4/wogdpuTGgoyZVzTQ
UGBExmCwAynHh9KoRHohCO+YIIAA/zs0XqUcCGq01MGZKzbdII2yT/+udsU2tKdHWZjw0PrCkOA4
LxQmgd8ZJB8mEb2pl8FSUZBEPxgBQ17QRmwmuswG4wnWkhI/K+us/+SABq/exZ/d1V+OkCQ87jHN
CY6L5xFiYTAzgBxYo4zpo+0NhH79fqyPP+8HiSdgsi2ABYjJ/PqBNoZ/fKi2cI7ZUqj/mmeVPBeq
t8Js1ckUXKVynLWhLpIp5LJp/wJ3S3bmPt4XnxzDLk1jjl8PqR7lGwAhYpVnOzIaMyqE4/PpqNM5
RLvC5xuMDk62RQu6O3jReteyA9H0qjmg5uRLjd01zQQ+Zs+ig53AQRyEnHXdTq+Xx2L2lK+p0i7H
yy+ieo06brwSORAwJAIY17rKukv1UtWgfj+Bud82/t/2coB2psCSWcCCUFPnCt8q+Dviq3uEEUbE
RXhv/alNO2XJpm80eBsrY+ehc5HUWQleISLXWVAQUn55mk3QFFBOJsecQ0qTixhGcwPiIAxjgqaw
mbaFScCy0gFgcyzRsREygk3C+vOBm/Cej0jyyY89WQk7IuRn53QRPM/PNP5uRXLzYFviaOMcnrmC
NtC0TIST4NI6LDIicZ9wWqjJM4LdruzhAQO3OmkV28SBuD3JnZ2B9Q+zK95YeZ448XD22LaNOw1q
CoOx2K57rYOz5elv2UwBtLnUVl6ET+pnGzSog+A5VRED7FbBNeWj06niTNrOPLqslHBh93pZVuzn
rPXrpDE1Pzu6BYMd3I8gCJSBNEnP9xkQTVLZBkTwAYtQHOXbDgvd8pG1wQ9rAgMxh2EOrOh2bFqE
+gUrwpenwjKK/4Fvk+jkq4V+ENX3IczeYI0KMumBMjfobcblZd9caBRfi1mwV/zgNiL4pv2CRWRh
RYyyuYJHWPpxtLNCyeAxdIkOf4qajtF8OEumRP6MEBDLB/tXtMss+NRVT2rZ3t9wpU9vMuEzBOgr
Mmj2mT5VNZHEMoXAsOUz4cvarSJOI6D7NIdwANVC7UNoTIfmtiJXdptPdhrCmkc4FOe9X7zmj1sX
PAbYMhEhLofbSxVuGdU82Wz9TaDHDBkkOc0MH5o326+EcMdTSWnk0ec2aWYWZX38YkHR1lHtWHFn
NNfqQQjX96Dy6nrd4Q+SHSb5OJXMFCXvwVEc0eHz9WT6xIiTP6JDioExbUH2O13PLl9uDg1W9Mxi
JEPXsSGl0H5vM9BnBdTpiHb1GTM8mj3AsLpgJDs8RgoSgiM3LljCrGIZ7JOG0zdc5ygF9C0Jgw2q
gm1GUthnsXP3ULacBOB2s6Q3qXeCPVYGv6bCgpkkXK57e4STqUHvW1SrLt+7T5F+HpyVwh4m6NBz
yCxfXEHgsMkZaNVrSgNFd0X4fk7M6B/HbJfBjBujq0Q+m1IegfuVborLexzgy1V+z792qDxJaZ4H
H3TObP1j7XbSFsfjba+g1kC+0CZgpIdJt0YUiv5lOnviWi1oyWXK8405APL2UUQ7etgHcT2yvvUK
kczzzjjkBilCIcuTmWHIG3OVx/fv49HCJRzoHyVkTruB6FYa7dKcque3Ss7hf6Dk4C7X4simiSia
Gk/8g5pi91DcZXWV2PxAuGaVk4LhSX4meXArceXGDj6gjMrhMN7YCCEUZbHpCKs60Pw1gyzfhtPz
/9cWFupm6p5lNSgm+SgW1xqp9GzzjCkE62T9zWhV3fHGqoKIhvhF1N12ilYs6LY55uRWIcyTsjTo
UaT/2+uvS2zpNmlusGCI8xh3WKK3ZWWFn4Ku8jeC0BEBUG4Fem7HrQnt9XorPHh59ayyOR4aIEna
eCtEkP1dUoKsdSY3+G52za/XvrEzcbyMzSql04fzGiTB6LFuXbqskWrW8pJJ3kk6AlXh4vfv8G5J
Ym6U+wDyrdNHcApYvOXCBXi1le0knItfL8lpLo/2xJpHCB0LU0zivJigE3GuX/sLy32LCMAYlWmY
8OSFPkBGIi7EiZZyHz4wgUATcp2SYO1xYu4oIt4/7jndkJ92M1rOLjnmw5NpqxH256cu97qzuYHk
my7c2NdD1Dwb1Ju1UF4zh0GYNBhxJxDvFLZMVx+yuicJweeewsGmmvdPxCSv2Fo8Kzrs5MVVoB7N
qKs2fyHV32OO0eHAjEyzWEkfS1RCV9IvkAyaeQWQdLfPLSsBSCTlBgUO65OAPLgcluVWkvnRb71i
B6ACNnMTkbs+42jbMoUei1I+2/7dtc5lrK77GOakjMH9mxhs9OOZQPxbhEI1GLryMY60LgAWpodY
y4cHumVuWAxgX1/+1IRTfpRjLIahZvFd5cSM5ziBHFgYW+qstABtXv6hXn+S/IlcheWL1OSrfQZ3
PptevlPulsT885zm8F2hhlSwn5iXHfi2KJMiE4MD2EIFeCAQA/8ktquKvsheHRG6d3EJty3lTLsE
8fiKrWFFOCN6dBR3rGSK4nWWzVhZ7BSh+67WQPKOOLz5RG+/1UTHR+E8tTXUGl7sjsAJDdVO+ZKK
wil0Ep7lunxUPBWEmKCARjb/LjnF3aM7+7AgsiQe0aAC0m/Yu2Bhu1LDxztWxAz7rAH0ODrw5R+f
e/nbvHmpYXLd4b2fp7Vc9pj+arGTwK5DQzSNdIVKxbm6HxqBWqHrFT+XVRVPCRnJIh4i2tT2gVXU
61bOH7WvGcMEbTIazr7YHArIMfcBmU5lmzsCdpvUYo/SP9QrvFLtEOLcmcdwX+LlXUH0jS07O5Li
L21WE/WPYyjUV8a0BTPYXjM+H90Eu5bdhTB1lD0h1FFOO73y+TFOq1kt1qetlvLw4M444J/L84sq
NzgjQjTsdKFl3kgPVlE/yyzD18bJdOq5jD9rCY8F/TVe9pZsW7XiQFrd9/1rh1DDB5Ja+GvbYKA2
4eifrchMty6DnPmo7sZrRmLN/UUQu/WNmrDLdi+D36gVKfzld0jxEZ8uAFdQDg1r/+qnR9tlyGY6
nE7sa74xHtoOMaoHqSYse2HARdGsAL9WrzTizKnuUPHywdjQy9KgEDhxyeR8O3rlLGhFBCIXsTgI
xOtSPD3uOXl9iViZIY4iYj/dhzYJp8ZZJ9WtUQPfimU6yhIzXspoDH9oO+A57wK8E+r5Ne6aJr4X
J8+0/iRICE1Twx682zty93t2yTzxznFV9ESsVvx9UQCtpThAKSChNCwIQYBJHngcpQyPtSFjWrPP
Zo4gTu1NMRrwTJLzU0QfX39alMteOvFEKWQaGtEUx3XuPxH/lWEXY8Fa1TrjpJ4Nq6EinubvqjIs
uw5ek24t0Hk7JTyyegFk/bndcfmnXKiH+dM742xv/TBbdZLSOL47mURxtUxn9BaA4nkV2xmXiXwc
yg9CzGwYN32rtWVlYVRF7URSqMBp/xOlbosZ/yjgRz5emf42BT6rdMp+p5HSLhWggHNoryKUczr4
eGQ15CRRCy+d81IZGu+NFdLbGsNK29shvEWIi76rFOPcul/UecIsUpHwdnz3PYjxFWW6G69EoG9n
7KHZf57pCyEC/ii7CG1x6a5axwq73yQVzK84h0zi1tD09E6VrpC5x1tmxb81vKIQpO7lW/QS26iu
+KEiPxsEK4unkDXa+BIxRqSUqvnckDNP3FlJAr8vema4Eddq9MvwZ5+P4exrur9fJHtoJPKRQVn/
ZmpeMPoSUeb2hEVurThQkGit2PijAlCV7S9l+33tZaXvNcznsgjISDUbknhZ307J55TA7oektCT3
VqBzw2wTOE4eTmT0iI5ToE6BDYViWUfesrkSg56XT34HkeTzWdm1ezC7zB+YQOAiihYWq2KExfU0
ONn7KyPeflSlT/B5hhQHSJCeAuB/0SN/qTSqeE00ho9Y6knQ8To3pRHHGhSsrWimZj6huuK+m+lX
8RJ59qb8V18qlWQZvR/zkufn+X5geqsQfwM5BicZxjX+8YlYi2jyiX2343bLAjv6WqSu9a3R5uMx
o2NvKxcts8x+oxGVm4Mo1WZQMecn0qzwkD+MbJ9FUkwfToEA6Hca8tPuEm1Io51WvEGwdCVlMEPa
DmvjKZx/+1k1M5e5OJXG7Mhq2oMX5QjCDibmxgv4IPqi+NOiC+I3+PdlD6Xkhxm0gg0BRPT/m13/
0GA5KXVKIzg/1/vK5tVSfdeghB8wnmoiXH7M4FTctlPlJ/wN+QfJz3923ex6Sdnauk+qIxOelAQG
B0TpuYUjaM/rNy5nLeQtEK08RyAbSiGqQCTOiOqyDmJNHvAAfsJtLe4kSpZ+C5BSsq9tPbZInviE
tcp1mfVGnr5xHnnjhtUG1hK4i2UB6S3KfSH2mtVsbZvWwmvnJQ+OiiHCwv94X7BhqikM/r4s5xDJ
yLDSkvpcNicHwtRgiPl2TDFNQNbg+mTvBbKiwKQxggh9AmFPTjWH35wshMDP8EfdNXLyW3yLNycI
QmC5uoZS4tOMZ7q8amt61mKU6fTsNyXsdBEfdc7URFQ1WxZ6U1WL3ekMr32IczUjL/KLqF2oiOlu
gfKEf4An1zVeu4n8RMBCrwrMnxAkhjKKxcgxWkBIqM8Ajo6VPP49OJ6xfStoAwGYSCfmdbQQGycw
HI1zf9FWb1kPunq+Yz2I8f0dyock8vAx51ClwwQ2IBqkHq7A4MvSRM/sVre7lpUV23x9NAT2x4D1
bziNvgPuK0CyMjyMYQYqgM85d2TMM9kGF/PYtV5TFnFp6F5Ku957hD4g71vgNicNH7YVW6tOXF7f
dt/fhkETWO8+eoECiNWIAc86n/8ipUoAbO+VD1EHwMVBlw7brdhRL1xRMJkw/Ody+DfJyGTLqD/p
/gneb4LDm7SBSHTjcKC/nYxg/Jmhx4BZZrCfHON/LVqejWaaANteHgpw0TmHGc6dD8eyrM/cX/bz
9j+9O4ul191blCJg/tsm7qO+UlgE7dTOGzIsaDZVAbuU3aJeyH/wTMdByQtbtZJmd82goX/ARwLk
wQkBNXZsz9naidmhzyy+OEcxde8VdzMniKdYuNlf+T+M6B8nDLDxbB6vz2heifx9GK+771PaLRIV
e0V/m00e2pKAhIvUHy/2Ui+SZ5HL6VuIbOccUf6ltnSCxgupLt0NzrYtX86GMpmlXJrZIj5TrCIM
ZcFOrYmDEauxvLrm2feAnxzz22wEMbjRFwAQQiJApygSnskSaxUbWphzre7Kjl1GXP/T/QZBV9Pc
hhRP0dccApWkK3htzKLRXcvl3dckIlqb1KgzCbTzRZCg4upAi9NUXJZ69zJsxu1aMQVSa0PbOONO
LuRjIVx+XRdxZO+36Y3EmTCvLGfUEz5BGG6Z3dCakItia7W75bosuKfhJbSYn6M+JAkv/shSy+Jk
HQaEMMg8QL1HbYaEia4x4WBOBgXhX+TnUDg5VAQPw+arxaU64ZGWYcqx/XoGRdyCP2idjHm0lcwO
/I2Vyj1cm/096/oSBghpYCwUi5e+uP/V77Skbe6x+BYsHiNZVEwVNYtm9mxzO1BWizECPouj6l21
vVhF4CaP3vM8FitG2BF7YZolKv0PPUQ4miHebvfrgUuXODIWGhejIMK4z27vSr3XzPBJ4jn/nSY7
qSGNrvTWLV6jppt9d8RBiUC67EFGSPodOTg4Gnm2bzTZklZzqh6ypvfj8LWdvetiffa8t908Ko0J
1nV1HO5XhxyrtQ67dg4yDQ2lNgG8fKHUbjbF5QuQMZhepyEXrlElt2MslXYDwXoEgqkb8EgCOk1R
nnfOS0MPj8Zw0akNcsmagA0Vc4bZQSA0hIFPDq8oMrZ3NAv4LKku8Fo1vsZz1DesNkxAWQY9lTEC
89N+ckPH2EU3iAw3qqU2U91bak2Xk254tUKebS20FwmRyevGmZzEy+EiWoTQW4pqnvSYFWptGL3B
RId55WIqtNfkgsSjeMV4GwLrqNtrNQnDNQpROu7hbJfLJBCHoMZe0mGQgkuvIXjs1xkMCTz36zlG
3t6zLnFEXC7gi3M88U+Jj871mTr/398pwM5Jac/166n/ecxnObojIalPjTkPUNbEO+tBYQyEtEpZ
jabMSh74nHo1+03kFQVBy/kOsGa4zalc2lDpd1+vg6gLhxOrgQxVsHG+Wxw4oqKtPF1AgUI4WPe+
hH21uu/NNrWYx5gqw7ACNWKKsKQwJmqtVsbgQsQKDTBROb6YI45adP+M33FsGC0zzJ6nY517DVHM
TwDzV334EZFJDjB9b8uq8ozrWTSRwBWyBFzB6O8CDYxK3R8jl1LV/cZGgXCTAID3eCbd3jNIz2v/
j+nqiDKXeL+AOJQvunQhqQ8ewSg8GhcdwnlFlsm7CVvON4wkhr378OQW7b+VuQTWt2pzBzXzyL9e
6xa/g6qxjkc7j2hMfquUZaHKse6hTOBbboP63alHvu8G41x4B1rOprUfbvmT2YvYZ1yyNEwKXDLT
bZeLxY2d6DRQNZq1ndxF/x/yz3XpmfGpkap15WDNf1z8JILnX7pwh5n54cZm5XjQ6iJBG8+wsMGD
efjsFJhyZ2E0UTLN+90uSLtUPko9JnsVguxxr0jA6jrP17Y5NCy8Ij5D1PrbOzy1tlWKFYCPYk9U
oslejMEFXCNQXLKk5Fl7W42mf1LS2qwOSbeqq3EoUhNdA4wYl2v8jG7OAiF5ufx10xskAoHcOqCj
GNwZ1qFaQQUZCKtYvhxioS5KnHcTdpkMBTmb/o3pOwq54C0lH62avovbkokMiK6xD4agIqB5ZiWJ
+rF5mP/quiQoeLMr4wOX0XrvTtNqxrw1Mjm53iWcpVGnX/3RWWoZGMS96iwPcwTxA62MAcywJA39
hJ3LfUYirUSp805zZY46/dApaZFrxVq0tU9ZVFpOQrXOTJN+xBPyGTIL2yRoa7yB/wg1VjmFnR8S
76R5tIZcz8uDaSBVMLx4ueyyABo8cT2GwXCAMQdJ351Kzn0nGH7a4UTX+9SR6t4ysE5hXTScGYVN
CmP0SX3Hx2oa/+ClRi4AdzTrtIBdLsEo0DSsmDHXNpidzcBGEj4IE23pUwVA8nJXItmNuU2jQK7d
vnUXVEEiBRqJ7iHZWNStYaRGaloiqG7t3putSt46xvxADwWiakGiawd9pKpjnM0R6UKH49tmqXTE
9Va4sNJctW4xmTWjq49XZ69n5K+8ASXz8ezUc2a9/+WDrxQm7rYI+b8nerujnD7xwSiaVzOdKnSI
U7dHNc3miaX7IknoKRdTq7B+d1dAVJgya4SOzYFlWUeVZDkGiEScsL5l2//cIIOjODd6rzYwt50d
5tmh9zMn/uSkfiq+Q/Lhj6esPJGp8aj6yL5/ylSqad2wKzgjSZ0QAAQbdP/wJ7n6ZjO4oiByEZ6B
ItqTWnwLs10b8qW6HmMrFuCCASAipP87MG81RX6MuWv5ygEEKfhq2LDgv/7BPBfFu7sJf8vQWbIU
KSYjy4tZaKHqZHWF0hVD4ewjZGUs4zK6MEREMGj876q8RCYdPcCb20mdf3/g69OcNx7zQP/p31ae
D0oIPHfSTq1s6eBmPjRrmoaDftR6k3+5wbWmmLllCAWR8ANgdW+ru70PDSf/DJ63e2L+dSuTqHuO
Vh0SVgwcXecZ3b0ljRCyXZJGV5eAa0EThS/Sih4JjwzxJ0XihMV+DwOdh7kftJzvuE1pgZ8Ah7CO
dFm1uzmIJoO5QnHDbHwfEUo8mvj1sTxTw+NkqXoocvpUmxwdnKM9vM2p1fKXQlkZmi+yvVc+fGq7
osmXS1Q9us56AVZsi89py+ccBRLSC6VHabbOj29xfE9+FbDgMp02U3W2sMypdG+iBhKMKOK89eNX
sywP6N52tmjytBSvzXz/kGcIpdy4XUJ2dAfUI2CWEqAl+6nCzwusrQx89Jet+75D+AR21isswOAU
2rwXsjBQlcKMJvyAbtV8KacGRh11sF4iUQrjKkOjgvYtakdLlCbwMpAi/nDzi4FOCgIvcBNSU5bO
18v6I0iKcUWiNKDUIfqjlQ8jxSx5yE8P4HxxbSKUKC40AC5yq/3XwPQjTXDd3ZDpvzCv0lwvQuM2
altyLcw35Nlk8/HSxVy9veVNnaKhyZm0S+F/Owe2FLvfg8XgVRcA3Hs66zVAa3t8V9q8pGxuRqKF
KbzfOJmvASAmpmFaamDii6dxwO2brpk1jm3443rqVh3wunid4OPe/O6JEXL1Gkfr+doe/AcDIEXp
rQ/k9g5sxP8YlxfR2Ck81IhbMkGM2UYZWLU9Umt7TpO5p+qu3Ncfw5RArjg2yQlAQULh5IaNJBJl
vik8kHtjlhrOny685A/fClSEnkp043c4eDMbynn3I+fuLs/AosMxVpOGBGf7gOaKyCGIttvPzcBp
I0xr7crR/4F+w7DFRcrBNtJuw7HHrcBhhP39yc8jtrhjiBhLwKpPABkVF1uRSXGLLZNWKdHh0Xxd
6eVNgOUGj9rMlQHXAqkK9XY8RXgGmuffEtEzyRHE88FUBIcfc/JWI8LRR3eZYsCyCaXq8eEomRtk
9X4jO+n4KzbDNolO0hC3P0Qu/OivqlDwHN/QD9AvbtFv8A4WxZdkFd2EkvvtQFhYvSdm23qdaE22
Nd805UWuoOzvN5kKcOgMOFNXSWVXVLZeA+jkvoHhj8Uqp1rR0yAtGkKSPkG/T+ELmYChq6gu7j2x
mFFyxUFaUMeYqkxBzhR0dI4o+Lu+F02JbUM9aZESXxI07jPmCZ+c3nOIY+psBNBAxWrKGE2WmRJc
NL5HIT2o4heIEYeR4JUsT+BrfeQbq87+kY1eD/MrfxoWRV4BefIiLBgM6S+Iu0giSlPcI3wsssVK
+JVigUtGCyrWFfZqwhxTo6iDeCrdnJHbVTyimX+m271jNKD8AAfWxyZVZsQt9nQKAt6kFmfMskzm
P2d9AF0SduIH2TW32bEjT+riqKSltk+Nndt61BzCmC4dlrnwP43GK/uczn7YCubZ1cK2kXN6U7HK
i1NX19PquL3YWdxbWKAw0MxGVSdz6JaCzq/Fv/0YWRm3xd/iMYnUfytWxQ/wwPAj38rYhx8Ob1Vh
pVLrb76+8Gn3VRHwLPUnHWg3lan7hfpdryFdMUhKNpWWqoPGt3+52M1qsH3X6dFvvS0OR1c/ALgX
PY+JV6UeXRZ9n/G0upy/pZbOQBs+rgenkL9OVnXZdKIBdGwMR4cKaXZr764sJkl6uciujKlgIrO/
m+0oPChTWDaLDNWwSo+V2dY7W5gw7m7ewfC3mWwYy8a/J7+u9AMY+dV5wDsMhIbbj5ZCffadW34o
koMu5EjchYj/+KX39BG1lTr0wLhknBOe9WTpcyRkkSqaInEXrqPBqsCUxd2RN1lST8kgL8Y+mtNO
/Jx5u6YuNCVV3Wg9396Fe1y4TO2Nov6TpoZM72sO8gJzpJP6m9pA1QrJ2JNqMDhoLoGN7sgHSOoM
hlzDSuetVlWk6TAg+4J2nTt0kN21Dw/eyEKTdba7tgb1xg0K8gBrjdLNslSHjO9yGFICuE9RgkP3
N/YGQ4Iw+TsXVLZ0FpYaLu6XZe/dTad2k98ajKKQGsDNukYKfzq8cSpKpeHc58K9WP5i3tBzcIGn
XSzFqj4dw2xBSjelUBtJJYiTfR7MVZkURyq+UrSuSjh8YGJapLV2crRtGxxoU77U8Nv9mHJt39/n
YE/lW4te0gI65Y4iQVRpK2Ad/jUw2QUYNXIIzz6UasBTogX2Zm/9vN6Uy/mDYswMZd0Iaoya4gPM
1FQKcW6joSkbR8YrKN0mI2oDpcGkOTR/04ESNBHPWwpTM9aAeKbME7jfSEWW2jv8ihsTJ3631nZx
/HpWdqM92DOOAdJJIjk1iwIE9CAZOBm1jCmaeIIjR3+a+Z6M8CVJyLXEmaCSC609BjDVw8Ff5BCo
PfvD4gd70zaluZKBxww8OipXMhcvqDWPAhBSq9aBxTkq0QzlOnNtPwkb8U0RDQHr78cN6mjGj9Dz
Y5slHwvVL8UWuEklhKKU6FKlPkPwnfrfpdx/xzEj++YwulAZXYMqy4LzKrsQyLAhOw7tP8+p4qWi
u+w6oPx4ggcCYSw2KL5Sg0LvYYXo7TxvixCGG2dj6pIUUURw3D6GP81qu79elq1BWqHyMzt3ZU9Y
EZdDM4/XgumrTP+cgO/H1Yh4xWS0k+P5YIFe0U+Oj7V7gZulRKpkdItn2YtWufO7G37d4zkOoTqT
tBpM4iLvLKudIh9jTKH+ksH0lGu62tCP3yhfZ14lxzsG6rbtirUkSHgTAnebI6g+CxPom91TEjSL
Viz8gqvp4svb8614CGhIHraWloLDkZ6fxq2mJm7K5BA285SqptvS4hMiaODW8ElL0BaNrlW37B2M
HdvS8mcsQBU2buKXi0yTit2mxz8IoDH8bY37SWzyoDYVIfjX+GMXU8jC+t8eJPXDcvnIYzlgYuFO
f8VNYBE51S/hlqxYmDpPBvNd8A/oZ9gh7Dc2/mBFPqxHROVDazpPyXHwZgk6rvX+AJBSLg8/wSDR
bSoHoAaNutCFuBBfmc1xuRXeO+gnalNWfnlhc3nGJSC3k6q8MBhXg+EA3ixtdtYu+/9hr/ReoAnn
caQLeQrUjYH/Bf/6MsNo/k8OzCiQifjt/UpY7U+7mXb5OGa41a+N+xwTWpAbyNtOdO+H0de2uu/s
nKlOl4HKLoy9yG1f2cOcTTyAI3DlIh5UZVsjhWEb4CUcAh69zYt/yDfnrKj9J1YXZhSTLApwE/nE
8prRUMwmtccm0oqbuF4+XnA+151kzz1soMyNZqLRBpj9FdZB/LKjox+y1PMaK7nRcnnNaMgxhHJF
wvugA+Dijc1aIPMMyISQp9GsCOup1qHTR40e7sa+p3ZmVpQIwWELLgfTxCJMc6iOUVfPD+PKPvOR
bEjialmxfF8kY0PzX+G2Q+L5l3qlDbtZWh43L5Y3TSOMU7xo05Gox3r2utYkCbdIBufPHq0i+0Pk
6je8UBm+Kkl4prLKGR2EQvMziyt7G50wsTwXO4yDJzG+n+5Khyn1j1w41s6Ji3KBumVpO5kEmBc+
moqTWsT576SWktj3ZyzXBzGOHlEAUeQL6fOWgoRtrjB32P8GWdtmBTS7FAQ9q77rsSAJ7LooBLNV
AFloSf1OZE3/diRWEwG6DY+AFt1+g4nevIT7beysGfFSxx/cHS+K1Pl8Z1QnU65A1zTHSUrbgcO/
yxlZ3pqdK7zhWj0aRwsD5ygJKcc2ZDoqdNtXWYacXoiFkrIsEMBz6XsSjee4GT5xqX+Hp0j8DzIi
5cezSPFST+nrzsZspFmsH9aM0I0U8iipK0V21eKpgTbgqbhJ4SJpst+/qXewASh6gGHu9yYEDcKJ
Xm3P4S5R9If2ZrbKC7to9zgd9qKTR8daDYsJstMDb1K5ZoYZrVdSZuZ+IOtOkGSOV4NN4gax0GOd
WMoD26mAji5BrynRf8KRdWe9fHIbd1Dh8mCpqhjZu/9ruWeFOFb7dsbf9bYACKbbj/SWiSUOaUrq
wjlKLKqCgkct2nJNZqLn/9HycMh1zQWqqtRdULAKPyY+lpXMXZc0Oea9ma8TZoar0dCU08BLWDQ8
7doT5P2IOlVHzc6+fknk6wFY7T2UFRuQ6WYQKDo1oDQ4sDbPXALOhFDAYdGemli/Ig1BdOOebIqp
1ZwFfVTSqxTB0n35XMFCoLYeBJ6Q/WgzYjW1e9rVQvlUWVtgnT11dEPQBhRzRTV4PXNGszJ0x0kX
7ZvJxTab4Q4i1VlmoPzoK6p3mdDGxCJFIi+vFTWtdWImTwWpzQr8ypZkviyg35YxjAxfBr1XCVtg
BbcdW4r+am2YRIZQVoFtH+B6HK90mNESl60NYFDsD5bCKstHGDnxJtFzdZyZoXwZh517O8Um58IN
X1thLmu6ZJHce0YMZ19Olq4hJR2IM9dPKzz6H5AmQHBIrGWetM4AmZ0H4D7+X9cG/fU+FgVNWhRM
6deZnNJy2pJY2sylaykqANqbOJHDT5f3kUHZvvUiM+dsft04vwwHrkHBKsMW5SuK8KspcpNdhpD8
rtHbuViPP2jaC/voB3F+q0mCNIzp4Odnog9Xl2UMSfcABXmdHhqY8VNkDxyWrSYUiOwiufewFL/Y
J2SPGtgp6ZpA1UzG8NwolIE5o2ltrxmz67SLjfpfNkoQn9/SgTK/lYiRW5rrJ/1oqhGQh999l5dm
hJiaHsnkC9kGstUMcBSossBVC2Z3vquQoeIyDSa7L9zm9dzk2OBcY8yo++2uvGkOX022bVqRQmh7
KA/F+a4WMt7+E5ObiIVfmgC7NVMICiOw0+KvhDRqYpFccGAg3KCbiezjU/J6P6xseVVYjTpmjqQj
tTmp6iUsr4OV8QZry8X4xLaYXkn3XNaG9OHbiQY89pi2J/ggN8jdbDQrfSgbrhPEJ/fzwKAXGu+r
UkXT/qMxGhQseKNV3RYRLm29WhY5R1XxGJbz6vWF0BKT1TuCi267QPEdNbbruMMed9TGF1x4R2Ad
NYGqXTZL2N9Ul0dNWRb6SBjwhO/m012tVg7BVPuTqFY5x0MJ56OQ6VIAR8ZdTdaYRtIQmGGmalHZ
ebzhlCyDZEoRUxmig/xeo5AWU+vgrpCFj895swKsHuqlos6gc4aQWAIl6bbD5x+np5HdO6hfTAoD
iRW3jAfie2P0R1GmHdp/EU0H88wStRlA7mp62RENr2XEcV0rjJP08Vfm84axALmWEtLwFwWjakW8
V3M2wHrifFJSm63JsUEXyCAILbxbfhvX+0kf6Z+C3qM2OET66LjgiqHFzIUs8LQkL15eaxi8vEUL
WJD1IeEYcP4d/uQ7mqFnVyYMWqzIp2X/Lmr7YNeSivFb98qtDYkq6b+aVYtQ7vqNx8xtZls4UxMp
+QJ60K1IZkyHG2uvbyiewF6l4nool/hloKln6FhV0cyEvOZuQPBYLyzy2sJhBd0BYgVqbKBNIxzr
vvUfj6b+zdWUfFGTZoVS2fDl5mpnMNEbkYVmsolIMRIkSAzcxTBgN8ZJlipCIsErkvXL1dR0585d
UsWxzmA6AB7SVpA0YP0R/fRtdP7c4e4tSOO1XOz8mHcPiF6AyvzTY6cVETXWuqEi0/cO7yEHwu8Y
kS3ToN2L2S10BXrQtm90M5mZ7XaOQpw4t/HJ8h+sEhYCxjMRmO71Jvgp8tUPcCbsFmXua9Q24ZJy
A5sBhmRdWEIy0J8RJTVodXLCAzESG4Qpa4IPj2XehCIakjBgSrdVyebOFSOX0+32VWQwO6pO2nkE
oX5pn9GEyvErpHON3TBxYiUf+NhCE3FUzBirBDJ2X7zCtcfwhDmys3pyMz4hRDhyJHyAO0G6iiau
+PESHuGEJ9poSB4aOPQFTNiPFvxz3ZeCPEVvlCLssMIzXl+de24iM9BXLGmhWcOG1Xz8gtEyYNro
ISUlGfFWvID2Cl/rtjhwmp1bnCQqcxNd/KJVMVCnsn4DFznjHza7vsrG4UZ5ju3dqG6cNNrYgAdr
QmohEJujWHR0Jt8JxoyU5h8NwvLWWtQH3J4z/XSHX3xv+r8x1NNQQbHYUCUV6xLF8I47Ncr4P0eT
EVkft0XQ6ugI0KD8hQuihfnroD2Y34V+Z8VL5mQkrtbR6Na9VNJuWEzptsjZP5iWDqyxuM5K0IDZ
rmkWVsfPi2yVfzU32j2UXvvgf5avjB30GwqZnQ2objLakD/tH2PP56IvSWBr7g2L6ZUpOJ4zhXeX
l8n8+rG6Qub0ier2donflrkP51byUk6Ur3Qt55/5z6U2zU4tqDD23StT0K1hwDb4QvxhyYt7bA7W
VFZykArReWo/Ac3X7fyIi3jbwWdDRaudkXSFDZRxelebBH9K8bDKCrsZ1txzfTImaseL9o3SboB3
6op0V6i4SvOhcndYI6e6u5O6+2f0Yd4JXRczRk5zK8SpoZiLlC7VhMi3cFwOGLXXUJ+mbUIAr2oI
GnqypfOogrJ0Uqb74bkTLdWvK8Mt76MP32670pR/1by4Of7PLFcpy63JMo330gZ6A8IqwRozS3R9
dPoNN8mDbyPH+3aXaCT2TTkgrrnv4mpZ+bmpxm/dEiCBSNtpSTvA8biLbWF6iqgK+ihIfHbHZJGJ
aMFdoGb4IP0aAsU/2d/oVUEaDXM9kIgQG0kooofOD2jE2TubBHYAifKiU93K1VuOVXAcsCD9Cmzw
RFEs0xBMH71OWC9my0JewlRPejGjEepAmiR0RysJwOEvVusiRG2/D/2+aM5qASPgBbahAUBPMBII
ZgeTCDPcYK6Jog0garauSxL0YP7aZP18vNS1zJE61Dc/2XUp0NJqpee0OehhXpmgL2fkjfhSqtUO
K0URSiSWDwxpPfcqGQya6wnoSThU9Y+b5ZMANNLQ9WSnAglus353y3FeB60Gt+sLfQdQILvr9OHi
dOqHzB0cnvLaOLmhKrAu8J8J436fEmFUFgwbiWKG22BYeSBsQ0ujoGcjX4zf7CQCJvGciih52Ybq
bvAlrKqAZMs7FA0OdYsrx9EPzgPscsNYBJs8TMBagdvSoAjuYU4G35C4Coiq/zF9yg8XeLRPE40w
Hy3Yz19ei/svmOYAjRiGswDvBM9Fm01AA8icmzcy2jUn/lzJkXSaKj95qC2wpdSaerH5W1gnw5cy
STDczU5Gawu0dm2Ja1LcqsmgIPMaVbt6dxymGtesa68tJHa7Fdp9dsyYNUKfvm4KRApWCF6f5cdM
yeUl0huDpEpQ2BVac1bx7di1f4XXC+jcj/pT0kqeBLmJeDi1w1/+ZBfxJglTXQ/FrKLwRZVe9aA6
4AS8wsdJtH+Vh7X1LZAyj1OK6DRRZQ0QDpp9eMgOHNnvu7DN6gjFyVWPJfMCGd/BUB3XCHCaGywE
iF9B9r+kBU2JhQr5LiAEiViPIcpCPjS0XoTq1SlG4ji8IauY8dXDDcxnhIOEsKbrIFt/F1m1PgYd
HW0B3z4+y49zE2wN5I+DJ2mcDPMjfvk09PT4kwySA7wgkHp5tkzM/ORKJXK+BrN3EHXFDx3Anouv
ZcD98F6J+KU37d/ou9EB6M7nfS6o9Ubz6m/4Z3drV6xLQV3Ul/ykxBPVqTbodm9TsbfWpdRd9nwv
w0lwNpiIn3Pj3pxv4Wcvjb0syCZGDrzNUA45PLptfrS2yNGoqLUOI502+ERaycomSOKYAtn8yK+c
AM8Se8zNu04rshuBi3vJ3X1iiS3gv1i+iC+FNeSf0BOBejqFeOhiSGiXXRyqch3yn9UM+/Fxu45v
Xrr86nXN8Ma4583Sy58LiSeL/N94/yzaqQ7oWjw1NBICxPWZU04+jPDqQRYybmofNKjwZhSdA3gg
PsWrQJm3UjOT7P5nSP2Rd6iwtyz2Y/aHbEhlXcYTx6/e92USbgjCsvK26blo0ZRXRSpLVflBVICv
Pi9pUQlb3cal0FJZLctbYenQ+u20G9IQq5aA4+pk+ZQQeHXd+/cZbWBL8sBL4wzAWt8QMDO3yPQv
GqTNbda/sj5nu3y4Rah9mTpZzr9wIISvItNOSumllU4WfGXE+XLZMWFEOhQC/cnxFxmYctj144OO
IMr4SHlm2/RCaZXj/vyaoaUBwqkzZWEkKNtrTL060xXHds5oilbkErslU8V83s7tQDe5a64xnPRl
iUCGLbGOnENUJjP+O4BflPjUMgCNufccDzDlSiDuAivpnFX5dZT5qzRYvufAdqFe6RnICCaDBfbp
nqzk+x98QhH1g9uoyl5m7H5MnathwWCb/6xJDfr2Hftq2SnPmcI2tmbtxGZV5ImrOVxS+tbOvrSB
ZFT1YorPvGqbUppJU3UJsTWFStdU5JBNH5crocCYPaAjM0lLn8t2DhRLruXFKISbMtogLJMn6tjL
/9upRoh8LgejjIEEGXxYJ+fPpps/ajplmrIEUX7TxLyOuvl35DbSulxBdKt9rOOkwWZILf27QNUR
A1bQDSdzCBMB8wJtzCQuPkqzcJJo5zwpN/3IiVy176Y6qejmIGhwapDui2m2B7jwm3Ed6kc1rGyD
1L4MEGGS/VTjEhV8/RfQQVfSJD36rh2f478cwQf3TcBJoU5uHqW0YfxABEr09vYHWns25JbeixHF
dO3kYvD86OYwdyX55Z/y0nyZvwgkImozSDR06blR54qgW/vbJLAlxS5/QqZ4p54J6kqLLqe7aIWf
WnZHckrgfmG+WaFF39EueqUGehwGdVl9dUnD+hq8aW8TZuxzB+gnbAlwVVL3TdZl6Sj077MG/6f/
1wzeY0UT7V3VZ1DkjUubJ4sBZOnyOCr8HVK99YHJrv+zGIvQe550zxmrbCkrHglw3gUdw2vo4VBU
P4bmoV0pHF6UndroKy7QmWog8pk57HZqvY5MOlWiuA/GarqkbCzyzWm3utIGi4s9gObwg5KeJk0q
zaWtkbL2eSrvR2TpW2YDHFD7qHPBpXtntrOGbwTkm6NSn9y8/vF9HeTHfFK26wBBc+GnG+WZqOk6
yqNjNAmZvxJNx8FnsRLw1OmRrz0ceMzzaC3oyNlxicx+3iJCtCttruQbWh2LndmvwX5/1JccbqcK
LRUzZ2Urw4hQJBHP0df7wTcI0difG2Fypy2Ex4Zv/iALdc93R1bx3eJddHzvEEbgF9bnAnpKUpNU
vmmBL0Y47e8dMc6kPS8XOhQiGjFYq2G1wqGmNuFjGz3aqK8kC+FWYkn4gOYQL7zO4VBatjF16BrV
V8VUfpwoTwWWFhz6esgkH86ONv7vGwFm0NrfE6WJRg42VAfbTpNPsQ7bKKaARJkIULIFz1zSGytn
59EPFWx0LLYaWX7v6ozSiJitZrGL/77HGLkcAMESFk6SXxhTsflEOxBfktLPgJpKuuePVWewUdzd
XSKaOJHMrSm60EuFc0F1azAuFzD8rZXDgLPVd8zPnl39AlUAvhPtN0i2BkBBQAfeoecChMKF4noq
wM9wgmAfc32Kr/7KkxqBH0BBxVKZg8RSFKfp7pr5oWfGOmoAxnmr453bn8305iItwHr5hKGkg4Af
itXjz3NZGkBRMCQ0eUZxzsadH+ktVYxmWG9FiUycl5w1/thErZEwEfCDo8bAyHDshwbRJcDOx2LW
LuE5RwlcnznS+5OC1TRbGWNlfEqmssvBqpkqFY5lqD1u2Qot+AStCP3j+Ys/hYz8iSyZZ65wa4QC
PoR0bFacMBHNMF1RwoMW0ExGgKF9vonrDYA9ZMAwAUNrYrvVaD8q+2gDEm4bcE2apUJGPkbA6LJ9
UIqW0LDo+MI2Cre2Df49/UfJ1Jm4sutFxMKHtMB9C3VPpD4ElVzvzlupapTcPJrPjKPV0mOlt9fp
OwjEPi51h1uFAwH62/MTz9BE2mtTPkDxJgmr3Obli1dn9q4yIzmfCVpmsqmFXpjNIlNgRCBgY3KA
6ABGQtxSrsHO0/DYe63bpTWqxODTTuqkQgW7p1BZ9CmhUg2yrl8A5pH/q7dFL7QTpErymzL/jhlF
LNHg/ZW+5ryuGoHPS78bDvFIqmi1xwXS+AO7gHweXfgyBJ7KqSehjPiIJlZYqg5xYtMLDmyKgY6R
rbnuSmvMoV+msV6mc+EpWLdzQZAk6yPIeFYoXdm7hW+Kjj7B2Eeb686HXi7OVkV4hjyFBhr5T5O3
5LCQlA+krUBdhnheIoVQZBIe5htI92i4S1MggcLpBslNezUnSLqlX0a5Iqtiq9m2XrTGYoVCBksZ
1pboT7B+ZNFZDGtkRpWqlmbQS2uRGXoNjiXrKI9MuKqrrjIyawWPEndpu87LoX+chvBAmIW114D3
OEwySOnJOplK0dkPlACGyG7n5BHyhFP8pCtZY5SRgpxUFuVZx770HYSzY32epWZC8guK6Rf3w8aZ
5mPHKOBAowTVu+HPtEaYcyE9qjeDEUTHSx9nhAXXkZZKgAOCmBkV66qTckWAH7JA4DIZ1sFOo0kD
zkSENnXjZPFtFXcm3xnxm71ei8d1rU2d9Phjt7owCJBlbDdV5vOwOWXYQw8Hfokzgcbj/mWjFjDC
mhTSA97U1EcObAaAU9uZe9Hli2TrtWuPj/Fu3OKXPNXRbd3HSr2nTu0KYYnea9+WiWgLX9NkkXT4
7NBO2xkr5Vxqyak9M7i14B85qHh36wBP+sTBtRH5mOROeS5dao3fkSqJ+yuhnGD++qLotFGjHKVw
mXI25Sdueh6/fHsLBwnQUGWT9SzxoSqvWtqmBER8HAwrJudhcbr14L9ZK3V4V/0gdYsnBKuszb/W
4bfozx4h+Zb5iQXUV7Ueq95AjztwgGSxnZo+gZCHG2JR2YWNrBotM6PsZjHihmPJXezThCSNWZrX
xRiuuEwz6EKtPz/2LIzaxBIfGUBxuFn6060zL8QcpZ5r9FG9NcwbjtgYxZbcbgH9d2d1ifyGKatW
957ESy82D0PkFag8hWoXy12I6Si3TvYJ8zJs+U7qiLxKZ8wfbhn8uUQz4pWUxK2xpyOblwyko1Z8
gyTnGL2CzhTnDesp9oQ6SstQaJJE8Q/qfG+QbbcYRvxX4cNt/Ol73LkShGVwElvKduAVfrw/if2t
eKm0eMXgXnsGgMqJnjUiR2O4aUl1C2MX+ESje45VGwRP
`protect end_protected
