`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XP4XoIQK6j5bfsy6ceq1KZEWN56NXJG/Ns3BF3aF5LZBbpoU28RGman8yEuTY6JI
Tb+hFCUTaQ7YFuARdRjsYJIP1cx2iNrkB8fZyCfrAOjdsUvxv6qFtxH1Mhk0aTAk
SidNeVF9BMN66H+NHDoEM26sMz1zN2avKtsskaSOmdg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11200)
FRZV8d3HEnV1Ygy0ZixgceE8b4Uxo2gpvrJxP/TZChjRFoJfwsC0smvc5Y/WnaqP
B2H9sjTMV+g9BbvmUgwOmGzl3hwilXdqpYpcSWPMzEk/oc+2Z7T18wTp6ceijMoR
TRg6alNeERoUFqWzcCKQpBhhN8rAZUExlP7aoNbJxQPDp2hPWicy5TpzAD0pKy6/
jG6zk9pX74aMm0IscoC+RaVwAI2T149rzF6ClMRst4/RWBGDb5gRfN3brg1Ka9HS
I3mPbpI8mCEWgMGNa+gyKQEyCRPSyWtOvkycVUO1K6a/oN+VHa+UzTdeFS09x5A4
0xumYFrMOiBngaFYIc/egZYPSDiXyLsrWapGNGP9uIPyzL6IxKMeACWrDv+Talzb
3vaMdjc93C/OMyELOk4YQZiL9xRdigQRh6KG4okZsJSL2iKF0a2R30pfHnmZlQID
aMi8T//Rwkx0D88IUGgxm6ScsFOFpElrWpkwlo9xWWAWAq1++DQgRO/zjSWbNEH0
NMxEC66l3fsyjM/FhZSwCNxNEIFoARd3Onx+2GSJ+NlMdP5E1enLWTSMtn9/5rDD
pPrJj4Of9X+WrFHJ5bOieolPsBOQGucQSQta3X0941cICWT4iXsU7LOB3l2sKk01
0PQPoFHjxKVy5eaW07tuC0dkmdWAEy0F9MbRO3yUXdYRXDyeCtycGu4UoqY47FKQ
ncQRx5dg/UwI8hTrj2fGc86nq34MGz11KuvoaRlKikUjXWQUJv9j1YA/B94QV4gw
V3udt8/NpdlBblpfBv1AXW/XsPhsM96k1qLcu9ry5VOZKiycPj9C4hA95sgYyXT+
wVIsIJJIJSj4/GPWAXGi0sWM2btsiPafDnIry0KCyxzf/RW/nmyz5l6+05zXUkrc
7+uea76mhhcKyBQZwuJEAih1UMOBvVZYtViYaVZFuOwcNJ3M1zBlYxl/eRqDCOTR
h79W83SMwUWCOjL2sBEhIS9OlT3WRVG7qnWN7V7wXt6bNHJFgk9wfCvpKfNp98kk
hPcS6iFhCTkoMt+jb1hb608V5X++a4ck3hbvTT7I2qT+L6LEVmBnEykKLaNBQYYJ
Z6bW6/2aoTi+AYt1uf7YkRAwWgcpKMqyO3RsEzE4JUvZIkoAN79mClOY4vX/Jp38
boVviBxJ8moHf4mkE1G2UPzrw9GHSlDIpCdG7/b6nRokyA52oH3TmwH08BAjstIq
14BmqjIAoU4HCHvjTLQkce+Hj23iX9bfBRYSjZlw138lSMwMGzVFVI+QET0LfqcE
lgFmcOqbyYq55HxZrhRZiMmBrHX9BR3RvlwhQOZmUzj9Uh7r8gOF78XFT6teh9QH
a2uEAx8AAi3vhOYmWxh/IMQwu7gqhtws4sd07LMbPjywlm/7ViFZ0rC93nXbyNkJ
1tRVqn3ODUZDjYiCHddepFW7RuIc6di4tfo5U9tJ4pRu2e+l6tG/r8Am5XjnxD1c
x5wpn9UWagSjOSRl0PV4ptdYuzscMx1qNrlunQ6NBrOP0q4PUdolb1EADIyi/Aiy
iuqhQBIyOb4BbycmXjEb2NLyTrQr/g36Yx3nyGS8wGW1EUERMmOxLLmjaxOk6vxL
s+LKw3oPjbd/ZoVYflJdt/t5hRB0qEgqjzsij149asrSYaSjdzHl4bLIuq9AQNVP
UlDd+XKTMJdcpdYdzehOOiPDDjz37iwpzNT6Y+frqCTIjTFXOxIpJOuoSIHo810H
+LT/NSJyq+eCa5CZKaMgOVvd+Sr5l2PfWQxSQ+jKY3OdA4CH5PAmJg0qozF7v2El
bYiXtvNWj7KLCh/SYAKhpn5I9l6jASTJxefX54dD6Gqcl1U41jd+lmsgfWkRLoVO
TxDgvWIZiU/jEnmtcdk7UzVqzndB1oqKbKbdpzhRZ9rzn5rDAOOGMysUYSC8dmh9
97kqFrndgy0x0yOU077pfDLqvn5ojNP2iMoearidXyULY1q4b/vcxQx9SL3dN7c2
syR1X1uCMynmC0j7bs96Wcuzx1SoriAkEOqJrZmmtbTI2lH7OKbJeB4IIKJxji3s
ym9uNVKxKNl8RMgQDBr5EfMPY3ucru04zbmc80mQWVuB1KXcifo8C9rlzT4q+OZv
a6/lyyE4E/NoUaNneGEeunMxtB/UfatpAG9Bm+MDrPVGoV9VOQtePJsECoHTx1Oe
0tvpBsD9X4koYojsETsJ7g5nh1oOtBmjGHosNLw1/0ltPPVvWymkJTzQ9AkTKeOC
IJyQ2r6/Xagm8hFM6XugbNUspq05Y0wdjQuJ1e6mw9WztmK0d63/fYL62bCZT8Eh
tTo+Y1MQuJiAqSXDlTUvCkb4KVAajUuokrCOV04tNyWhKUuJiNZNOTQV2vj4+CSC
zZv1pg+45wVcJ8R2Loet/qBsb9RUfsJMz0np8ohRrIhqIOlSMqYg7SfjjV+NUWPr
UADqyc1NIUQH7Xe5d94qQ7C8M+p9C4BiW7l3WiKLiHkRwcEFR7PgBMZVED0cP9Yz
IQDByxsaCRYxgWpnFHKbmafBkwY8CWwsMcCz6dJgQB1jmySAWI+ASGREKD67qqE6
28MwxFnZcX+aPGStAtUbw9B53RYikQgmSWg0QE3I7ig7/VUqHN/ZuBwifNkcp87y
6baobBZytvlMu6x5zeHeq7HeTlUmg9UCDyYh2L+w247uArMoGIKzCaoaEd9UkPTo
9qTuVEDQr8FlJs8xlkpMyTN7sJbPzaEyTp6aS8VwCcyRYQxr6YF6RVtq6FNIz4NW
t/V2ykyfzwAQ9PV3dLMTkyRJduaez53/CM3sV5qgF5ahXhDvAcoRM7ne5EeAAQkY
dO/Di57VggSyHvPIStXbKkWr4YYsjTyEJEkDi305KgRw8qrV7T9/lQMsjShE05ms
k/e3wkHZuKVTjFhQTT6Tm62bK6QYu40nfU48eY8D9OYPPfxGtqNUuMC6MgelSFO9
E3HUWstE4IqO1iBfoeRy+7vas5c1HFXfDNc7tNFYNe4+rZTLJCxIkETEMISrnMXZ
nls/k0s1zxa5QNIpmZfAU8aehuPDg/iWh4inZE6Tx8fIazjggSlWGkcuPZSaUrvQ
C3Zsc2Z+9JhP+hJBhSDDN5vtLTx+9fJILwCOh5xbLlpgr9crVgZpJ2MMAIk/kgDv
0ib0KQMIneWIyLfj7v+3IBmFXd625LUNi7v2+pKJWUPn5Vc/DARuBEYvYtuoUeTJ
niinMNDOoUnGLiA8MCar7xRPdc7gvwu7D0UorfDDd2ET7RxjMJ8itlqFEZwpl8Ik
4MfAqmSLW14IWw+PAg5DCmn+LFFC4o5/XsW5Ipqa3og9+en5vLkEqGWo8nyX1UK/
XcjgO47cVYP8auiFmHZ/fqXxa3nYjn9i7Vhq7cTf9ovfH8L5mjMjFqeUgZJqN/uf
na4LUg198IDupdSt7CALiJmg2TmBtHBv1UggAxVe0rMiAqD+2beqt5LzijvbuHbR
ZEHdgIHC0TFOlg93nOpAY0nNX0Jm29j37DLe5CREliEKV/HuPqAeaei7x48UrOt+
QD/PAXgQY/IT7CF51Wl8Eg9Kz3tss4BGEBQc67UWC4HXdE8jc0z0CfdPVr6NNF/b
DclJr1t/U4u9ddV4VvCEzGrfnQPfRflxbtVZFK2DSopbrPA9ls7QvXU15bl4YUwg
PqIgc27ynBkXpSJ5R1GRuTVpoV0Ijua3Ud/6Rh+y6eMvtpzSSsTy7ND1+BRChTcr
/q0rgjPKnN7ONUd4/MHgQ33edVth38W09STeKv7J62ZOvpzgiSitA8kwNICJSBeq
DYMfo0j77CSdn4eTGzG3w6UA4uKDf2jv4GpNCTZXV266sNL8heYSMdf9GJsMUXQ7
kk/hnkzDLzRdqmmBKBal4YhUM562/B52QGrSar+jgSfCytVLLWiAmt0DaBHRMtuW
Knrn0ofWLm/lBGy1C2X9gCXp/L9gxtIQHhxdqNPp46wze+eOx9Y5tLG6OWPPZMAK
w1Dr3twEwZfF6eOCANYZK41fn4XCTRvRJDhphK3wmm+4Turw/ffHv48BdMz9dHDK
5OXFI5jEOp/ArlQv+NdoWCM6v6yscypy90JbYFDjVFkDRogAXbVu6XG301vMbfXS
1UAvgBuo3d7ZIPzAGut9nsUqWpMWaVNZB4gHgUcY2JOUTRg+GKEdoXd9d82E0vFm
KjPLg+Kfy1Gs2RyMzZYlKjPf+xXZNyJUPEb2zAq0GJbppdtQ7v4vqtm3oe2k1KnF
fK6tf4P9l2HCmnkrPJ5ouerasxohALr9EnFdCygGd1Z7G9uTTjCxdXHbT4l/N24E
q2BOedSZBb4GH1GB1FAThdn7ejL0DNI9JucbcbYPHGvXt8DHEP0JikuI5kgj2cDt
QwXDdmlisN2h/gG0b2qazYgGV8V+aSrOjQdOA1GFTEoFfJBAcKISm/jonmI1FPj0
yt3KR3WmQTKoZbs3Fxp4fbf+y5wQM+GMnvtyMtTeKQES7eXA5tTLDzgMvrfWl+jd
MYya3cEchSiCpVzNyE621kG8JBM9V6XpdG4x+tglZa+SxPqmFnAuuG1VUkORto4L
Qtw2rBW40K1FNOojXiZKQxKj0dlLLcFTW8JdrA2VvW+mRbrm5+TTfHlv5pdcSMU/
4yvHsdI5lAGW3wrWH4/y3igSlCHrprALy0hCXRZBmewp7ENP0J51wa7Xq+ToTvbn
a0RWYEtOlaGSTWhxY7gBUg86TN88bBn6AcN0VywiWO7HbporWxgR18dQjBFMM1n7
Dri9vF03OQv7ez24/FQP9J8bawUEO1hG8VAfKa36VggiyRqZsAGWQYcfSgIYlFCf
E5NL5VM5hjQYIIcUAKvx6a/EERq5lqiCKtEtSgbnBLXJ/XuK/KdQt6PYq88VDme3
Tz706DfdxKjuqMbL6ky/IyZcDm7f+NGwklwfe/yYc5WIpmx3NSY8bsk1fWZVk6FB
grlQhQx5AYoi4JY9SrSyZ9lhnK6Ty4g0kY3m/ln176MTR3wcPKbOsx1zPt/0mR8o
kB0uVbkuukUW4vlC/iRqGLTA7kEHBJMSF16aJTfERbetm6zCz2O0kSfHUdZ9BsrL
Ilf6k38nkgidYxbnR/XADqFfOieTHemBO+6hTQ28XqwHTScfjT4VUxagTfiJH2In
bR7EDtq+Vc5s1FGo+ejSOFEc1orCdERhGVvMMAWuJrUF05jj+wwUOpH7xjHoSXyf
fN80nxlZLxF9v1Fubc6lZwtPCmy57BbalZ2MVvqiyxWhsiyVkKi6KA2N1FYFceJe
pwoeZNDTAmONroSDvtINUo3wtY13Tivvajv4z6W9PfsCyDUq+aE3tn7oTkR0Ikgq
LoHq8FApB0gI18veMhrJvw+9PObwapaQQ/BIF1QTQ34yaL52Qb+HwxZM0iOdfM8J
yN43ljkC7FHax7U9ZbqvQs9FkQaZOHfcb1FeHHYFaAiEUEKuC5jd+MjezJkdwGOS
ts7z7s0zLUJ8l/9z0gsI8KXPZwXI1a7znkU8tnjcOg1MFpsqig6Z1haNuA6ayw4z
PKrCXVbQc7fk3oR+7AI1JojewWXsjV30oalW28SeRSLwnYjmUPZdHCgssLgWXLK0
vKOzFopVgx+Kndu/xngOgpZXcHLp3bYXltvWPnjiAT5c90xllH5xUGRXpe3XWMTy
X2FbTJSxFdF95E6uLl7sBs25aNRIaNutgDaW2MH1KMX8D1ATNA4ecUV71a1GlR/b
tynn6Bkl6yoFzTh7nC14AfB8kYakev7sH0F/Higfht/8/nRNy79MPreHtQwpOvBV
gfZMNocplQBnXLA5NZXBIBmAo55wV9BesrQ1RCosy6AM9gtZ9BsoeP7AjLuD4Fww
SsXGaK5LA4aM5bzzxizq0reTCS68kvpVmWp+6Txl7WolqCs6rEyUv+TZT6b0chwS
1HhMxlB/Y287mzDDOt+suuTlhaSiyrw4OEvPxiMFiLRFiT0Tbp/CY5SDlv+Ek4Lf
znr1WuL1MoL3wlkPta0fY81PVW4bGLGj4PdcXLHbCFfyFlprAFX7nK+/CMazpiFb
3eV3jcg+tbOLVHpOcjj87l4NEmITHFd3kcQ5SytKqhz9GBzrooJ910UQHgJzwBnn
wP0JdSUM2eoVOv5xKhOXuKQpu5B6ZOzzRiQ1VdPPTVDmsCDp73iY3c79kjI/Li5a
GfiV4/tX1QUne0U9DaT62cftA6zjC8lqcTHW5Uv99QDwA5Lo344bahQpJ9pMj17N
gnZ1JIqyvF7hLs7EvEXd9ihHjygHMGHLw87zBQ4f50PbFBJx1dF6hQof/aP3sALn
Wz97ZW/d6fhYX6t4gtpxefdVfwwDFH+uuztP7KbWaDHCyBQA/0pCquNllQAf6PsA
QgMtMhwQlpWHzxUeRFICaBsHN8QSyYWdT6FzjUS5U6KULrnm6UFuzb8AqnWR/hH+
RNf3o0dUynLZhMZUXPqnQcrzfVnByU1xhAs2hUwmF9XIM5e+QlMJYZVwWzYzgB/k
U2vMCao0JxF+Ivx1ACn3TZUjBLN7jHgMFkfDiYkl0bNaTHUNaz+4qzIB6pAL2aQp
qJGVXHxzCd2S8OEG4voTdVGD5wycJAKHehEpIk+KU4YigspA8roYphkGJ2erdDt0
Lon2ngiU1V8EsscLXKk0Atvkz2zPnaCnQz46qDPtvy1UbL3nU41rI6JE+hWYZ05k
2V821R9l7KIxL/dnIyZeT6UjNWXm6zmBw6vRIvGOrDqsxR+6hi61s1SwVzw+FTOz
AXKiQRrWVmpL4g22nb7ngNlGBWUbXIVvQ5OaV5Ygi03EHiy7VBEK/fvSrsWxDJDi
zVv39/hGsQ29Jr/Yf2HU/jdKAn7UuvwRCrFKnkxeOZeL4la3bOI6OJaircJGuPWB
b0XSlOyj7DMjxfvX7GN9VadXwsLHFrbygplC95Z82BGZHyDiB28vrrbngCWKoMGl
lAsdn/o+6jgtx9Ua68bdWWMtfcwJZs+y0E5Vdw2wo0oBwba0es8P+1kntOVxgETB
Bz4BK4d1v/jBODNl+r7k/6aCNKc3dNVaLRfkz5EbPTYsX8pI7QG4B4/EuB7dfebj
jpZRnesLoHaGDyp4su9wr6XRySO8F7h4jWby8NWtrv+jHLEVvuOEs7mFCfLQN8UQ
iwOJj6OZ/EHoB1W795e/pWGUY7k4UH3uqAXZyBdzxoI4w/AiqG++trtCYN4/CITw
NCmSdJxi9c/Z2aORR4ehMVu8J/Qb76AdjNyOBaNqNCPXb3nGcdEiJv9ZvdHPLfFd
xOeNgoc0FhAqWN0sfS4ZcZ3zdfpfTcwoXy/H0PJM1tiOH2+B/ubrqYnleIZY12FW
t+oIQ2d3dhuEM+zsibhR0hA7EDtDi9tcZLyDdnQFXIYC2T5e1m84VIMlyvNlM7W4
shg/gYWw2I/QNdclrNwlHWZ3mwGWpEzZlKQhb0C08WYJ8He9LtT78zcRKE5n0L9n
xyHrmUyTJVwJsvbkWJPkiU2siZiuZAKwxFj6elw93XIBCIC+M1q0EvG4ehOZr47N
bOkJdGOq/AM5jl8Ojpn8rjDcRw0KLXGtGEscJ4Qf/9Bqnq6O1Mj39PMyfKkD8RhZ
Z23GJzYebQ+0tOPYh5yyzhLP3NQanCKn9y3dewqYyTrsn+0N9J94H+m/6l560iOI
JgIJoyD9fW5FZG0jp5tY7UqHDK8KenJjX+uh4+8uf4rkRICU0S+dfpk2D3ygFmxR
R2H1Kc/32pGXifR3NJup+Vrqh7ELh/jfSEM9CaJBsgQ9yN/JRZmxQDJ8wRWnDJjG
5svmxj9WYttIlTGpgEbBS5ucEqSppJA5IBIdXEoLauokGVdKwnqbyGoLG9Bzgnxa
EweY/fnyFuuPw1pB7YjoYYCJh3vYGJ5XgQl3P9qzKpwaEHbSz5XPMlUAkV4H9B06
/9cAVEAnwUADiwC5b6/uoJaWBsHEm/p4ALui6fxVvvE1wQKj3qi5Po1eLT81b73f
U5AoWebHUfrUxiAJw5dAeUXMl+HBFamPa4fuIgOWmVZvIXpX1DUexgul2yldyNfr
q9XHvpjXeWPPGIzk8MU+xigDPsLbqmuQk97wrrxNersHL4lQgD4nHIML0EJ6g+ra
Frjr2db9pQbp7q4Cbu3TGTeCpv95fXZ7D0DhSDyHDKh9iFQMRLnyGnCwQX8zd0qw
Z0XMXq7Zr0WnFOaItP27+lu11g1ypO4xfPTNs3iGdOYDz2nyFM8w43QsVsa0GmE7
mZPl/evmk8zWA43ydpnYJW9hH/ebhHYOcHCkR5GJrA5deURNj+npVJzQ+8vz+t7F
tfVfrcvv5hoIT6dUh2mcZVMvlPwHyXs9G6O+55YkhOSLQAL6ff2YyG9tk+DQ6mzj
xaeYYMIcgjgX/6BXVWP05pLvaQ9Bo96OJ5G23s+EQwzjPV046cgsv2uJSXH1WFOb
cM9j8ceY9B04BJopHK39WHiuXcYHhcfbstUlufxVoZoTFiQ1Fk9vqK7rDLrmYyLn
PqoYLiInm4szbfgg2OMNpsVD2b6o+TdJxoss9qzxrC01/JYRzZZsALLgEuOnms6w
Ezzjs7aG/98hdHioNh4gc2/PaL9gL48aPvF2Me7pzY4eHludAJlu+3pkGZQW97Q1
orvzfONH0gSlItkBtKfJjzp5ZM+hmyNH4J39gCFmfxngoVlFMEJlg8n6BKVbeTkB
rvbsfZLPsFOVrg409TcRk8Kg1RvZSwd2UFz+G6SEks0oGxDhwb1RP2q+hNBT/u79
8nqR4WnDdJjVmgVqydrjXAmRmS8rbz/VK4tDzbtGrJWkNME3cZo4uLy5O5e8z/iF
yQQYHSU2v+yAjBmBU+OUeQfPI/xEmvnjWkPNeCQePvE3ag7vbLvFARBaqvG/i3Ps
0gSi12ObBcL9gzqIlnvBE9z0HOMMm7QiirbgfM6Op/4KNgilW4mkvXv19DiBhkp1
YdrSOkaaBFgMZlJb5XQgzJUfHJ5suyJknhbEjkUUGFIUGJ8tE403iA2IpkLPPWuL
ZSDZvnahlhJLeHOAcqmmHQusBDLCRApKS3Uj0Wi+koGJyt0PB5SzAPQWhxxh2TOK
Tmt55kl9RS7aBW2c4rYByzbEbbizoKbTvDY9jTNiufeHM2ggzfCte9OlQUtdfr2o
APUCAzoos9N6MdsbeSexnN72YKnuPGylvuO60RVfLICAdwapnP/qKA3TqB2k0eiY
L5TDA/lbVYfPtmEuYl5X4z9hCvErUxXpb0SzmLUcW7YaqDQvJcG2DZUJWBC+pe1R
ItcdCw3yV1O93ow9nvvKSUWGM9nzErszj+HfnVKRZuVstBSZxS15Undj8UBP+kiK
Kw5UJ5qhZT0ZSIdLVfaTqlc7MJnZGeyX3cO8jAJEGkXLKy/gicp9HB8svfyAe+bQ
IfNpZ6iPR2BDSciMuFTXu5BNVtVw4OQqu5PpJWUG3zIFxec7mUDZNycwxxiLb/nK
ZP701n8bYtX4rgnE57X5Qa/8mHMxLF3p5/2ycKNHNcdeHUQ759vYT5diynn6mDeb
21A2/+9IeT/7R6aFYn9IYselcpJS8XxJwUT3+KKZTa2D7/Ln4qU5seBG6jRE7IoQ
icdoaLAWPKh6QWTHAjznmzRNvd4HLerXhLWSFMGr8vWtPLYo+cndAw9B8endaQNo
vB2nX25Ke9La+/9YCHUBm+R1aPzFj8TPLCwTHudU13tIFc0o4pO67g/9wMrYAR4J
UaMFWrSODQ1xczOfKXULiUbWC8Aa7FrrIoynGbXJALuwcTfBwnsSuqEZ+YanlUkY
qMSRttAltv3uzQVk7r5HXYu7QVgiViARtVAWMpVvtUzIYBnCc7ErOW6l3sw7Q+Jh
9AXyuTllvnWXELa0orIXHAyWU1XDgM5gSaicoqYnygdMY9ryycfhuM0jC9+ykelF
s/qTeV4TVaN9habDlUN32D4JpBhWY65hdcI1i7SUIrq/yNWQfjdABrs0OsajD+Sf
0mL1uu1FAz6+PGpNfijVRbs8dbX7jD70N0XlrXo4jQcsoGH5f6sjT7bUUk7W96nw
lXh2ScjCNuevLtInK4yjT4XTgY4Dc8cZo41zy1B1ReTh7iRAmoqbtebP6+kRDxKJ
af4yxrLeFYGf/nOn2EeobAazo5R4PMp92CXOPZL0mdaoakoz4T61qktc3Wv/FKOZ
bIEMJP+skLOTozn3DmvpYJGdKmCvsyX5o5OKnpsq2MOvkflMWXLEG0a4gdZg31vV
HalZ3CV4QQ9kdYLcQ0NRdEVoeJ6j4U4n95+SC5z52H3gwH7cHxDEcIDxLGPKVw3T
NBMGfQCX0LRp8fQoXSfdZ42d/jDzPji297gnZy6H7MjUH4B67pKK3Z571Cawgf0S
v1djbvGtaEuvzt2oVvhsyuCF3XzwsxKYA1OVgkX6AjY63eJmqTIPyo1TColENZ/D
QwXVkO1v+wm/qp3o47d2LLoTPpXd74Hgq8cpIoF30ewbseKcSy607EyGHBPGZcmw
fMoWIxGMueWhj8tJLZLFM6AcqmnK69FmP/wGvAsAvCytFw39FmX9yQM9hrW8y3GA
7+7Z4ddM/cOv3DyZMTzcwI+xMLqyp8xEIoVe+3LVbmRsuRNRViTk3oy8qrniaIjz
sI0hwR48Oq3d7QEOz3PyT0g17Oviw6ApXml8mpL2k9VmOPOC/S637RKGJgQ/Y7xU
ACtHlSxguE4BotRFu4uANqjQJVSiaTym9mKCaVI+YKmtTJs7tw0CFk4EKMHx629v
e+jaB9Yvc/9qq5EoNwv0DXVykd9aVxJ5lbcYy51R4dQ8IbebC+z31GPXuhVeRGqE
ox5j/RoHBE8o9GchVVA2kyvxUUKlkaPLGPeDDToH8IAZkd7gqQdOh7G3ZGrigY2Z
PHRzjY1msmdaWeqLDsTJAUccqtKEHeTWCmTC0n/Otv93OLh397DxxPI9YilQ9cGT
+1wwBAOYw521mx6jkP9+Bz+2krrNQt0M2VwnhtpSb18YPPx1rD5YLns6+pDcHzQ6
dKcgc5sm0YW1eM8lxQNNx5R9JfC2lG5SnJJ9CZBaavfQVC0LxwpkfyQ6vC41tRDX
65NO885pG5OBSPpWG3c1pAvvaQUK00D+XjryaNYHCeN4rXMkricdMYF/LS210i7l
6XnvcwCSO9z67Nvojogx9dAWYyD08QJn6u32O7ivSBSv3uKDYZk2y5sE/x49sFz3
iacgIByCGfQUO0kJJwg65V+IbQYFK/AHfpp5Br6augaNyKN+C/j8Qe2CwM/D9l/V
X9M+mOSiPKCkj+jY7/l2vDmzrRGpg4RU4SFe1kpPjlJRPe4EowgLIAHSdcn0jCO5
o7y/ggWZ5ypF+cGZZPI0K2oEOPTjvtPHonA+BRAwE+YmXvRQm5ZZHadsX0TfS0u4
OZ5bJthVz9gLTEyBsob4x/gGNAHwQA94Q9IuoKPosJ+yr7AbBcBIoC/vTD63tEjp
KYETLkBUoNQgP57AkbVK6bP//xrCfEGfMJ0Gp8vpxRRuFY0jJcISd31d/Zs/ZrXu
cfQZi68+zfTCPJih1ehPzfvtaKwR/Og8mEiUKzXHBH1QLZLz8Xqp4ASLsd8kulKS
WDEC8iE5AUEKTRlWF6/VhO70WNQq4hiZ1QagsyxD7ZdsBKtqamvkHsE8MDs0oYnv
piG7G1zXh7H7fOcDJJjfLh6Q7QeeKY5XGL2GBnt6ltMIOhskpkcnWPu8TX+eGyRA
HArPe3f2BLhVNjqMbeCqaxFSKapuKzco+Cu2erCt5kFSKg+B0tyPpzXLy/NnMWPN
vFn52oG937ah7JOmLVrYzyWaBf220FjBnpKT2i7PeU1rs55NV2OX/ZfMuI8Kl1hV
bKJ6MIr9AQMB/m0fA8aBdJi5gi18X32197Dl5rdPK0uTSEygNdq6ISBhAi6OqZnk
/+A9at+RIlj3ZfpvaPZgjtu6EPy1l5ZbYVoBNm/UxeGkN546L/Io5g1V3yZk7Ghw
mA0/sQh5g9yrIfR58OzjjYgn+erB9k2BXUuNW5sz9aW+rVOyPbe9F4yy04rC7TDH
CqhWfAxGIaQI6FFjaP8NV4Vvho4TmAvRqgN986GOqrWJHpQCZfxSZZlF8AArgk0+
5JriRVuwfVnHtuQsZaPLio/XnOh0/rUQxtdPzv2E9JyXMj7xCcjtv7jnrOmKg7PP
yIrWImJY/GN8HsDAo5pYLDhEue8H/vVO9BwQFRWjC6oOS8PW8Ut/Of5hH0ONa+8s
KwvxZzoFtTrTP26CF7n4NCjM0OW2S/lgLafYuLVwJ50XTU+oIXzZuaxI8ArDnD8k
qwvZZe5e7hp5rflAg3RJjlJucOLyJm6MdDUGBs2lWD4ag9DK4siXuHAKP+NVD4Bt
yefRQwg+DWYhz+qSw5wqjkW+01xEff4AhE2OYH5b2BPPTBL1zW+8x5yk61FhaaEZ
A6TE8Yg9KbJx9DHtIWMEQbS69ALU3HBDnlGXlngfV7xhFpvaAeMhWFuEuDHWhQl8
GspW08lhUCjH9m8lTB7YHzKVTK+JE9XX/qy/2ra0hUwzro3OMk7nBbXHeEW1cGQc
KrnztazwnVgYDqaagU+ujbRxBBdTf6q40Yysa98yruwYTmmy2FZ0OwBnMby5DRbN
7YPnkkLjasm8ptQyIF/o0Z6PQHr1fLTFCvVuAVv/ICnkzKG54+lEIYXVmMzRJcBC
rw9nMoYaGqfUbWFLzYxjHM3WvWAv3ZAVOV66N5VDM7JFed0UOebVJ7GxZiDUre8W
WI4DL1cfRBRguqeDIjBco7o4jMJr3D6+xSConWXAtfJsgW1vm5OPmPJj4YyKMKT+
gFWP8LyilF8cO0FC5bwOBSNoWs6ZAH7zYqd/bycC2IY3a7POek+OnfRBKkqbhq+T
DHcy0ejH9uOTaN94BFmoOlMFUjlCXiPybMfn4CgFZY0UaSNHEG6ScFxZzBz7M/yB
xOr2eylg0Kup/JK0OoJ9pQq45InrsHlQ87OL+Do2L16ZvKETLf+7XIz8Jiccv4F6
CYAZUt9SFQakicwNL1wbZHBp6P6AUXF3KuTyfhaDgnVAucUjUg9y2HXwOEVrxg//
HUSELBSWtRWe2wZm8+XIpv2uvvQPgB8r3BQupY7r76HO6x7sXGlhzrPLqNzF/vp/
iXxhvrFSuDym6WPCm1EFkbHZrrVrWHruk4TXBXz7Mfg9U581njclnyAR7ZIrzA5Y
oocM0IDk+ynlXcNvihPZXKdVB3yU1lpaOigVHHs0bkBlxXVO+ebOLU0jbdFh6ELH
22Adrv5ZUg1a7eA6Xb3RLeOJcyVVXVXrNdCqRBvw7/wVub/TBKTX3axy8A85UHta
25LDiUaBvKoxjf8vFOrGIQMHBc8hpvYTsOUSYlpAjtzMxfcPYPmlUGAI9ZAFC2s+
8h0MKerFaUEE/1eaRT7JdZHV/G+2E+WfdLiqNMNbBrW+aYtnZCGPjT8dKRHS0zhj
+o8xgYuenymLzCJAN4pllG1+UkFKanpA28/nIG2Av09PQnUslfhwADIzfK/xBCP1
uR2K2bbj2uSEJ1ve5OIyU0ihgJIcdSzePS3U2YZH5RlIwrKFfj34ZBAP3BV0P9z+
AvNXfyc2/3SePfRyConM+J5eJgoMfarismhIMRDPBYV7+mJMktERJI6ZUSTZ6aC7
aX9NBqcVB7H36Imvqp77FWsRNGp3meVZrV0/IM63mSNZpa6LyNFLldIgIctu76Se
sDA+U1jvr1QHs44wnLtQH2wq/zIfQZ0dzomPjrGdiBuiwlBnjws8PpvnzkQUM6VG
hWE6e7jAjLAsr9HhVBur5LAYbjKw4H6avWjTjfRsSch+8G5t0DwK8kFE0FnWqShJ
47/4UCKUbUySS7qVMEso8EIr5DWVVd0jgOJP5/u2cCfNrIWOosUN2Gcpmlzmocjk
ak/C+mJSYER1hk2MMuwnUvZGzZyAwN0CzPbZoAsWOb/IiD4PkjxZ1dve1Xey32/0
zKik0T9ehgiQliHbOaYbOoysUXSPVngzMDOc3Gv40zlq1k2Uqs7RVRCj65wmOhwG
dBxU9l74a8TjeesZ3XoCTiFdh7icF2G7q6k2o2Sy1Be6TwK6We3worSP0PRL9ppc
iX8I+UeehGQuS+rlz+Fo5rchjRItPYcciVeF05PfMY/kbOxFfNKAJYEH7aRzo/+J
sHlhLY8zzXzxlDfGImRu0olXAT3/Vl3iHCEBagRvbUTWUshTvcE/DEmM/LrvGyji
45sDCdK2ABVqbYvXT279v20gADFpri2PFZE5Oh4eedl1zO+VXKrtsjhU4KHmiKkQ
4PHY+SptoK5RmUZITrM6R5/2qV82Jc2TQlOgwRSZzgaM6KItPY3fezVP892plnca
8eGAqUVtoU0sS30GCaOKrvbQwsslS+N7yQ3amWBTXE0SIZozYx26DRQKThi8hQFy
tnHVnKaBkYyZ8r+4yYCLIGL+GEm4hiGK7QQ/orrQNx+AQPFnLNYRxXd/UMyLmcAW
uaC/ANneICzs6YL0jUhS/6yXx60USsMtvIY97KTAo5N+7DseZKfosHwFa0MwRAIS
KvUebdOwfmldXspW+Jjlh7x9ULu640YLPcAcDC2NHiODcXmIwiyQKHQP0vbu/SZ3
NN8f1ofwxKxr5qz8JYwvyFAmxNUInR5+HgARylD0TEnUfQFaFDsxI8b+sZqBmstO
6n5AFFcjGmXFWR3zLe3QOXgRLdtcFo1Y8k1mTfjmdD5naweUxF+uo0I7HhxEqYn5
Ss6Ec9Zkgh3XsTktmMJUXVW+OcBq1L/DnLMEmLYgM3XrQZwYI8vgjqu7MvgU9gWl
J8iZ1CR6f+TEVuqlnTlHos91dfsCrJokvdrrGgYqgLWy7qKUH6ZTcgE0etN5Uqds
SapcU6mB3TDc5p8k/QcOPreOwg9kKxVNvIa1VWKwdyq2+JHpuTaUw5A690XnMJbA
k5IPK4UtNzhflD24PLi2T6Qs7mmLqnvKK59Q0jesqHN4zpWehm/oKNLCtJHnVyd4
BU0c/RFAkhvZNXU67vQqjA==
`pragma protect end_protected
