-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OU0s5Vw8UQOteNLFHDHpXFOPUz8KidM2IV2DszCXTnzSYuABVSNcTGdcXGOL9jbjoRzid40y/CyH
YbiSyO8Rdnj9czA1sotUQ8bo7CDtLkwpf/yTU4VD9DE5dmXuggUHKYK5J6Ln/B7eJJs4QYhQFBdK
GJeXkTXafyaMvzxJ9dh9hSaOzknjLk300Jr3yj6dHuyD1X1T3YKZA+njv9PDm6n2ys//iR75MvLb
/IP3nyFQG1rWr6RKyQdMMukxUNGtqWlUff5/q0QAxhCgJMBovKqC0TalemYwGW7vq+n+L69bH6gd
XVYHimO2V9kLNxdeaMr7uSLe15yYooBMe2SU3w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24704)
`protect data_block
WTKegOhY6uHE06u+3EyQvVBzuy8kRBnwxYMg3O1oPAPXj+78ZbzgVK0DWOCfpMXvkOi0nOgMD+Z7
bsPGtfR6CuKkD3bMaYR1RlE92KH0cpI9RzWcT6CiF5o13rlEg6HVeKyd6dSdvX/oOcCyRgmCCeP2
hvQr2JNDogSrkkNwfbbmvBTyg3paK8wkl+dFY/89+c6t3qCYCPfY4fc4pEqRBxkDg40SCxBhP3SB
A5p2rwnnLoQIxXTijoe6Nw3a7WwqjF7XCxNfKV+p5GzOLJlgQiOVL7Y1LYbIV5VqR2zH0E1JybQ0
L28gBeJFXqFm/imULwOBn4Ju1SyCqvx2KgEPT+ao0WdqBnA7WZo4IMYrln8Tb8FFjI9nAOH0rNS8
QUZLCedvLD/cJOD2Xz8YU9cmiH8BMVLb4mcGLVDKB1DlwxgWXmH4Og/ceDZ190ywxFSUYaKYl3EE
3hKX5JQqjVvCkq8GupXUOSBNf1v1t8yFtjKrTiViE+E6AmxD1hUpGakAspwxJcJfi2lPYByX2n3R
yqoKyqc2Vyd/7ASbPZ6aFX/ntucgPOKkHG03BOFZxAVjuKR0qgtIv2pqhqXD/lDHx8qGVIg/hVsp
o7G+vj+Gey1s+C0l4q0nShgSCdg7IMGC1zhU+VgLU2qTpr3y+WPbv8UPYMOyMY5/AABshrK8aN9N
EUt4BqnsEKaXm6bl+J9eGBFDNjejLGDZd6ks6EM59vpy4J1S5xjvDB4D8mIPWMEfdSavWVMrgD8d
N0rTiEXWt2OYu2sNi6fi+JMjxpsP/z0BTBfm4SJjFXQh9zol43Isx+F8s3kIyXxkvpZuIm+gwRxl
V7nkDwNc90aYEY1pRpE+RW5scLG1nulVTIUYTz+/z6hOYRb0TXgkmPKKv68fQkE7tMfOcnrCuHnZ
OcSRfOhsf2UqwtCr/ZN4Rs3tKlA9+quXGguYe2swoQhxxwhHYXKl49ZiEc5nnEVPW1wkTsIztNEy
p+XACwaYO/KvSgIHMLrdn3ojNlSeWravnjpbDsTVNq3aTt/eNcHIWLIJB8murn5pxtZ+GLOR1IlT
i/hh6IWbbFopdvmNU/ihFnzPUu2OEPLz52yOzkieGlWg3RUGGmm1YPM0nOThN+uxoZZXw5+mNv2B
x3o3t6XzoFjr7uFVUVPf+yf4nTU6d4grGtz+sRjFPVp94AMvlbSTiAPxTbp/f/nxxGFGmdhV3zUA
OaSExMSfFJgy8S9E+E55FRpnthvLm7/LNXRBDOPgX0YfO18e7DQtiVz+PZvLrfKH4faB4G0u/RT4
wU9lm3/T15j7lz+3ldfN+ypZ/XFn68uG3jNWVdKU/rsyRUEbSTV0shKSO0IWCZNiWP4hOSv78vj/
QiJdVR7Kg3HYt5g1yEhm0zGuxJ21cE39awJ6sjgvJn9buGx0e2K5C25f88qgkSrloUrGRffY9aVl
DiIbXXXTYC3Eglc/hQ2NxY4vN38uhPgoAoGAPiCCpYj7Kamra5r9/BZCEpcZmSYq2Wicrv7EAAY1
jP5EsUOvbCFZ/MgX4ekd8VtIZUXmVtdDDW6Qb1yoMXivn76rWLMqWYipjpq1Mr2WshZH/hir9u95
D+U3GHAHY5RELkRr8ewnjeY/xfCrK4y/PltRJBJvEvvELYHqiPWOlrwCkFE4EA65pkfqEAHyIcWX
MNyhnQzNI+WCaLb4ZL60xfRwEpFAc4coqocmaH/msSkprczGOJITkI+WYXthYB9r3B6DfvK5p0gm
c7H/hvEXJ9zfDc5FDLhtYMA0lvKHmaD7EHDFMYZ/rV6JDe8EijnDYqVTlcl4FNoFcksHxx9oSbLu
/2yrbseE0+dEYpYI7FwF+GoYnweu4o2kemmSTvwPR+dZOZFO0gig5xCFFwWdpQXKm0Sp57I1SIp+
0iRLTLxS9MtDGrOtHi698aRwo8yk+kY1EuvTkxCtTX2IH5sKCthfMjORYkPZoup0uQ1KJMqFY28t
m/gT83K/E3+/yCwUyPVtdGF2/9N6aPAgmePmej9/Uz1o8Yw9hdhkWtQ7e8DdwtQvKzxqFVH1p8vG
GAgLmk7PQS9Q2fRYWEc9tjhSw7yQe7N/++8gPQszt9UFUb1gClbZSkpYLdwQHEfqggZ/ujRpYG7B
KElAZI5ZG2xUvm5XrEGzPJK4A4B/l05fRYXyriIfhvMKPB7W2udE02j7oTVP9gif5ZRIad6eitza
Z711tBcIoRY5SXGZ0pL/g/d37YhyUBJX4Gl31wtz7yAFJDiU8/LQ0nTs8wFAj2vcGTLi9+sXLIEb
9WkzUdxrcGjLbGuvZCHmwMzOswOCAbOjPkNDF9Us3toKe4b+x4BUUXs+tlEWk5mz5gtlQ84gF0AX
kqrKU7VuRrqd/2/7SSGM/edsbvWYdyD4HpqctLzjTMNDL+ZdpzeJ42qTyR4mV9TpbKkdxLcnW66J
qAM5qzlzAthvb+8Vo2z9LBiLiHTBqrZdW6Lc0pkymv3hUgXH4vIAPyvga/tXTDhEmEJTX0mFEkQI
pIQQrchbxZkWOnPT3aOIf9kgdSJggSHHWakPZeND4WZhS1Lv79lQXDdGsu5w423QfpdmQCXhCrCJ
aBO9sz+NJ85CkFtuvFrWY/wMqzGRAU1aScmnqR603E+Jjzgc9E8Wfs36r86GL4yF0rtqb6ck7GRl
70hfd3p3BwoJ5i805E7cqoMbtKwP5GA5UbAL97DVrUwU+0nslU9KmBH1Cap/cU2icoYNbF32pjJA
NJ8tvS7ixO+wVEy+3hH99Uj59A8Ih1QeZN/t5c3BeX7G2oqxowrbIqk//ZCUaXND0x4EiUhlsoVW
0r3Dq+62ZoQw7p6z7+GfDwerhjGxPn59hQuTDtavV3SIM1REy67IAe3wcQ65BbXBahqfs+FJhnyr
o3AweJ30Trif7r1y1cqGBUcSUIxkV3JXoBMZIMGWC1C0jwJFQR6hzuoxdl8vzNOoEcsBNMygPCeX
pcedH8b1+kGaBqB8TF5DDCxuEwAeiP892NUYdGQe2buIG9A03Act50hKybB88Km6o/QE3vFBp/ax
W96aqZfCU/bUzqZRDdf/gf/Fb3HHYX7ChWf7iqQdGdkgWXDZEaRjTFhgFBg5oWe0BhImUJ62Kv8v
kqST8+fAIwzcLPRP/akxeqL+ns9TqnbTnTsIZnsAgF3p9gN1yV1Uhk9Y/gF9bMpP22ccBj0Qk4aN
RFXA+pxFhemUXTjQXy7A3Eek5aT1BwAn/QErNcP1JRMsLu7iBrQ+wiBPU8npAsM8zyGzpFeMRo2e
49SLsdZhVqMfUFtyNnrdAOhRjmOoHb57d3VPJlZRONzEn/kuE9Z7lVj4D7XqQ39T/hFdRR5/AgD3
XDBUVFeciiAmImnJf4XqEJDAplx2jUqGJr8ubBZndgULLJQDYevlzpIZXrsqO9EBS61vRNIwhbGS
H+8JY83ZGvzEc03KpiF1f5Z0jZH+Pnp1uVwEJMcCXo7azPbC/WK7PYDU8hvgxfwfYucMJIOrRZYw
1g5/UXk3U2tBnw+9jBDWdNvXLgCYAFutj3jcL56BXHqvR1Qu3E7szqVh3EeESzTXvh8ET/W9VI2q
weWUz6yf0Q8tSBpVCtaCs3ifze9oRFfUELdv4j/zXJCtJgBr5HgMzcTh1B2AJmlMaF80P7KeAC/G
8yWGpklKdEyvewqNwNvcFr3Q/ojNN6A96Sbmo/DZYc65Mgn8UrsMcM5RBpzpR1zZvY+AqBWOdqtH
5gC+o5+n/fwZj0Vue7mQRa2tWq4UMDAGTCez6Gg3YPQLcyf4alXvRYAMdjKWNNd1nUUER2qap9j0
JyB103UqEsHSHNo1EnbKQMxlhMFuoPtRYHF5Hjman04TEWmpbP8h9QRTAOcwCyjHV3b/hT53MQF5
tbaYjMWEi3utcZl4AlwljFCES3EEf9ZrRz+iYexd/GoTdfCsSybayJYiX/+fPvukJhrv/HZEN+ma
nSyVrytILZXwD3yS16WebDwC/LtqTA318IAFKEotcfYsb7nEm4nbFjbzrynHDzToqDwn4b+8UO5I
Nnpm4kzxPOhM8KNwC0JBSF267dszBxOvN1ULVw+eib4s2YZHOcMzpjTujtlOh2WmtYAUF1sVbJdt
ysSGfgQN3iXtSv8Bw8QHxUExGdqlSwCVHnPVTI9Wz0THp0rbjgLYcMxty1OsD9Lu3VRZTSFm0lcz
X/oNeaTpA3qc1Zmwey55Yrvhfab7XAe3f2eeNPq9346TJ6OSZrBb2REGGaF/WkssX/vnEHlBMV0+
iYepQFyEyVgfKQ3UCcm3J8gqHbeLZV+wDhPpV/Hj+Rrwu/oU8ADfewzomse4v8QARrDEMGE0DmRZ
u5ujCmC9JXbSIroMgyBXhy5K7f5ChJe+GqSwk4BncJUyLBrpUzdlcsR5P2K0mL25jpkYl9PZcfYr
9VpUzRwm5wGL4/XcfUschdc0M0Khxj4fNeOmgYw/qECUqAUI/G60hAPqI9p8/S+BRukA9IhqCDDN
p1JmzjB9MgNL+wdhrjmA1ZjfG8QSua+vpoAACLv80LMYJHBegEjryPjtx1YqbLaRpmlpdLhoQ7wY
XvGXffMzfRgvtCUt4BCQkr4nqmIpGuvBsJJK79jwkpnYlzuxmgSJZEBBocLNI5dBcUViuFM/M3OH
FgzhJANSAtXElvqD8jJvjNW0Nu4/t6hfeRhECmNfVcjcPhxC2GdHCStDuMZQfEucmxWbIyKQ3Gko
MnCfy+b4aiO5Fqc03KtSTY1nkvMGLGmt768ELGttFibjAqy5gsDGZs0Suvav0PyWan8MnLxhGSg1
7YG6P6+8g/vsXj4YxZEEMOXYbNiyCINrdvKW8J7Cmlgw4ssGrZvEFSc8+lw8YCMbJ2xU5XljIcYh
KH3zUEO483fELYZtQlwTRdyOVLT2nNeC2aKOE5XRMpXRwLcASjQq4LBf3NEGFyvha564Kypm2xXR
Fqn9V+LZr6/VYWZCOShHmGuCyyoyp9x54ivr+BB/SC5oMRQi1ittbR3r7yH/6uQk1gII1B4j+VsJ
1zZTFuV1+4WD1AGGlYIxmDv0Epr0eDL+Ahe+k+uU5hSoeybStjH4oCRB+2ihfwKc4tcCqVCPa3wr
aAqVka21eRrHlGHeDHWvsKTuLSB5HXWu1FHCnY1e4MzslvuNpk55nhnLeYM1gr8ewRxRoZNvjsbN
/eGsN5Z8rWj6mHwTYCgrX7PqUmyv5X4/J6eFpaGLr7adjGP9f7kf+R4EAHkVorbPdlHACaWi1Z/i
qcWd9FxrPV9+gYPtlXnmS3lLHQpW/POu5+Wt3qXjS/WS6wO1cPkc1eo6UJ/OvJXQR3w0YJiiTFEZ
H8Ja8TdRLq3oNov/Be/qRZjxGkI92p7M6PHTFCLI87uJAUgVFxmjxd45Bddo+cX9HczE03/mDJxc
HgKrTG9oiFgeuB3IG3TsKMeeWhfCO5ttWo0cM7WodC2LrIvQ+kxOEP/mo9I6ix3eFXaNgWyXgMUZ
s3VkYEN/Ywl3x95GiJ6NaSY9sN4xn227NOpYBElz/xTG7CCqVsxQ8GObob7iv2LvPEsM+T4hiCZW
Z8xU0BGETc0aO8eVgkOACM0WF3BJOHCvA9/hAO8iL27JgpdrksLFPIapvgdV7JQm5JdF6AT0PUpy
yZe1kXzSTQ2LBpvFUva7sdRmXq7amC/IYYlv+kE/1LoIJCgPn2BbnKKRlvgW2U8DeTuddYLvR9CG
s7CkR124bPED3SssVXBahAWWDc/iHbqcJ8nZ0IxydCZiaW6mGSWwlGkUU5N/gJLr0kiYte/MhqCG
yy2fWp5OcUs8sNYxRKaW6/PkaQnfDJ4TrSo0syUbq2UdH4V4gQxzG/9IxRMx/fa462FzaD1k87SR
8xk/X+ZksklO+vZBMnpLMP1kbMYB2XpmGErXQA+CH436h7krL3Y7lmyqCjELc4dhEY/5XtfjCXak
Yw55xi1C8D20+GEtO/xMXCNSrFVUkBqNENHU6DOfJuoAUtMKI5gfgdn/H6SIpD3PaupCa4pIiR8P
0W/GzRfPr1JEgE2HuG4qewRd82q8tbYh6Dw5iV9F3eMm2f7hsQlxXyGAUSG8CCS4gxnwUWh10jXT
nCPKmpYSFGvPAXDvxGb/mZnKYpIwARLEAAPXMhy/Y/7E+v0efU4bUwx0zSuThG6fam//847nxfQ3
2ZCkxNwm1ShdIUYZ3VGHSUrUVXvAugIyN+vSRCKzU3wieE42OgZbw515HnPCwAgzadr9vV3krpax
7wpAx2u6IUZ1n2T+a0McimejMxpmSHTz1ahjmuzCyMUXfASh1sGaPn0oA+dTYV3j2If7UcAjOg1m
q4GOhhUaZm+uwHCtshCOyk9Toamf0/eJA1wy2lqmnuLpie0SMECkMP9MI+hylqSKV3NaBzVFbccw
7s4r4m6d5tK4T8yrEvI9H6h+fmRSzzZWpG9Vjxp9qXxJb56jt4zwwzB/+hCOldvQWqoz0AcG8AsV
Aw6+gqGSLCIRCFEw1bLBdCogjdDI30hN1z3ibyO3YH0uSoe3TWFZIkVaF6KzVTuzAEzbzktd7Suv
VS3agW6ySU7mK87Cu52r2SFMBNVnZOJHXYohu1CID6JjQSjM/wSWn01zI8+UOOAcAZzRX4ypc4w8
wp2+g3H0hJYLsKtxo2Uj03bA128LyifkXrL7bNuDBlaoWj1fiaNtRYj19JDp+D85Qc3uAnuhKNLy
eD6gtprpJDejFuONY29OnVQGJC9iYdexqh79mI/4AHGh4K8/R1i2hDm1CoiYiGadAh1gH1j1O1K8
5KEUoGJjYigT2eglso4TCRAu8wpbLfsmO3nIHq7TCi69dNoM6vdY5Ja45TGC9cGuZkvK9N2s4Irt
I1S/0tOlyh6wiUd3e3JOoEgwqhAuYi6+dy+BehUlc8Jk9Tk5zhgf+ibo7BjZ7i4ZnDYuWL6OYB9M
lTnQaJsrH/B0ioM0dEO2dvAqSLhkIRJo7iPhUXKOJ9ia8KrNF8QGodvLSVmSpYFkp9pxvGJreGp6
Nf47nC0bq6C1dt+vgWxgG26nC0xMU63HPiojF5+oSzBsQ/vytQlHSN5RJVMgaSyleQoWyrKfrtwy
h3lMegUxvR85+bFgL4jko+NgUF1QXjqhWIVRy6+Bxn67ePh0F5W02f14quH6eLLgKnsOkR2LFqi3
kYNkvDHo5kTS+7aLEyQwGtHZ8QychVy9BjA93GixxaRlfKDfjGaK/D2nrCUroG31RMZx9W+dtsto
LKpJAuCzNTlkxwBFHBjWytncXZcLn3HiYeNBiijdkVgJdRUNG+2kcb1CHNKmszr+7iPmFKHwbFgo
9EiQVnN0/LqV898qdVhNLhAv/HIciyeYZRaHWjTIjpY3JgeUOriC7hN/50Z/x6Hb61fyj1PBEQdV
lujwZKlpznkGenzlUFhGrvDV2xn1ZUjfJ39oZNPK70Y+pAUFHmfJKdJwr2cdiJDvOYDLLNonFosV
DDvHzcRxh9tTep4vl1clVdUk7Y6x0S7g61XhlGe9ALGPdNj9B6zxkyXM8+Xbm8OlEUdBO/bbu5Ex
PDbLn6U3Ia5fy7hWMXuHnZXLiJrV0vCwofZ5tRKuCU1wl7kGTaasQRkGxe3+3Gv41l+EhhTzZol5
P+Q/xg+hf4Umg1Iel2lU5CLj5rYsDURndxSCmGiedFmRaBEi92ehcL6TJXGmoZ1r/1nT/oxhPwSQ
K/vI2KRUfnzpv7DbEAtLQ3EeDMzkh/h3vfTQmhqZ1Qc+yL0roh0ZnZkt/1osCsaC3QfEwlyBIoPR
BBH2fxBkV68DzqT3bxjaOEHWcPTeTgnCXr2WUKTfKLh0Qhhhos8cnLnm4aVPbPTnyShyRHEdRQaR
NwisfeUvOkBJilH+sVhY+lVmnuW6rrPDqzVQ8xAMdboWcWUwdiTKTumlSn4F/2fl+PRDZkFn8xK4
va0dW8Dj70cA1pwwKShlOef5WU3enKb3hgMviUcFs5ZgraJsNTipcB4YGez2xiEYh8LJz3FeddTY
Vv/4mk2LmtsOh0W7qT1XZ8kVozpPzvoPy4x0+hbs7OxpwMLNvuy9fuHF/T9+3dKNot71VoLOhXCv
N3zt/PVRf6zpPgTNiqx6txqxBJvVMcLYOVt8I4urxRbDGarRb/m23UWw2boz+niVJCKFstcASL9b
W+ob1OM3H/E5JynlzGrSvJCiPeKjFkNf44AVyBdPJAnbrxk3M3wuRFpwdg0YPiyCv5TrRKalD1IE
1ZtqydQqCQ0eBZQIhTbDRu+9ciCqOF0j97CcY/zxWFTXBxtQBMfFnYGfuBrKLuPzygQ5S0V6eyDW
TsajNjwcJwe+bsUensKmeZAdX9sYyI+/QFRPsR3XCWE26Nki0M73zsOM7FlfE8a2oH2gl4d5Cdij
yDupU71InEyMW2T92CMhlQZtFy1Hna74KxZOLumzl0zsr3N7QVaod7v9GiaRm0fGYmTjqgV2YvQ3
BOoJGNes59uz3Vc0Mygm5tb9gdL9fnq24XhXtWSs7mgJeCIA8j0L1l+uVSUrxDgtwD2I5c85k0yF
+4R4IZpXpUICEuk+UEqBhl6TWJAcHATTg5bHcK5MjdTrlTlaIojrBstr9Dd80BmjIlGECpxXW3/2
0zjpEZqfpGSkQzskX1i2TR/SNLEq9JH5pY2VuRE+Wbu0FwOGWnbyA3ZqXuZOQ9+rM46sS/hD/lTL
C6zqmDLdtsYtriIunSN0pkr65gpX55mSasNO/63KBXLByDy9lRVHSgEwaPK+74oAW2pu7Yle1QJV
CLuJ2N21oonsCCJw5v6KAGJ42KmnBeideDXRYuRfPQ5lHKGy8nBmwJZo+d5gb0qyp4vHsL67GYwo
g3lb3aZOnUrR12GzGqKMfEWl9rGWDfCDxRN+A4d4q0GVOQgQkGfK+qx6l7QS4jswOV9z0DEYr+Ar
HomheJ1okwfTGtd4AJ0SfoXhJHrHwLWj5To0788TUaYRRbiBHM1VYjre5oWaF9OECXTmJwEmgxEx
T3Qj6bvbPE4MnN19oAzvntP4NddYt/PYP3yA6E2e49+c/UXM75ad3vUxNNNSBRstA1/z93iDQWcB
5556GYAdi9laYUr0VogZDFEetLLl4LdgT0nTZQ3QlI/onKP0MNxcu08t5aZXn3BEK1nmr5gVxn49
4LjXLsy5jlskIQ/xn0/KEejn2WU8v7U0/CV2JOQvsxOUQakd+2Vu6t+mFATJ7jRvQBbO1FEBgxPF
xrk6W7UMB+0z84ETA1WOkE7Sl+BP3cucBDI/CzODFijmpm2WAYzJTrh7doutFsHMWfRWILLHOI76
9jJM4n5Dt6UNNpe/kdEYM7Fbkc73KvOFcKhW4bQomMNlArtCJ2Lorsm67689LHcemnkPDxrcqdC6
95jrZijyQx+0w5mSaKj5ZJHC5tfEQ4MMOQRiH9WUtqxrApXJgv0aQM1gm9hCuLsbSzT0cSoccG1g
Y+Dam+bhyCDAOMuI9Sd1eVnFixT/wcGHd4dT7O+5AK8LzAxfjFO9J99Ji02SFZtj1FELXjI6CcDW
4l3Jq536gFnwqiRoG1wthYq8cVBZ1S6h385Qwcnl7lG2IPTM0VgxI9uxBiNLJN/SSt6HfpTghuvc
CDnZQewd78XmxAmxUfbMt55jnrG7z7mY94hpme5smMfy8ZTr93YLjQf3RdpDNW4Vc28SIoloV4bH
SqIuOM8VZ+c2smHuoWTf7v1WySr7XeEPY0M51xjJnJ8H5gVRy429y6sc3FMqYNUihPKFKtaAPsm7
rEEs5fqAYxmYi5Fyk0rNpzF4F6L4BjYYNPkjocWjOzYSCBt/2kHl8yxWbSrBpHp2gaSmC+JUxc+N
I5pPt9Kc/xBH5sr2SQqYYrJtzxVhd8opjr0k6ZaGC+Xvm77R2zYXCj8jcX4z3AtiacCmIwAzXbYo
XTV9PnMKa5d7Qd1Dh1SKqyU9Ddi/Bo3cQDf49kUMD9TCq6Zt/JDrJtwl0fkV1Jzk4RaRUlgXACJm
iFX2eM91NNb4ob4t8RFB9x8HrlFYIuu7UOVN3c/4HptbkYs3bKskjvWs4ypO4+frPBxIll+Cnemn
vM14Nf8qdkPyL7GxOM7i2zv5RS9pcroOKswf0MeqCRoOr5Ji6B+C0Vu2/Ksmne3f4A+dovcq1Dut
dtR0W8ju1Qng4xqLQOuxJsdwveB+hgw4SUSs1jP+OGZqsri1f0wu6iRX5jyc9L/LBqSAlc9pZFwD
N6LogRFg/C7n1x4nWhH4y2DhQvU3GG7jMVXxMmc6hi7eOa5tIKL9uGR8qrPbfKLNXjZV3mjc6IQD
ikj5JeMLtziGx6/E8+XyaHNHFMr5CPvIJjnId/1Hm/lFdLXF/VdzRfCNTH0Un8xGocE+WgVjIpI3
gCz7B8oFZkIHP0Va89eH/Vhq1GoWl+qU9U7T9X0tYdVoNnJMgk9h4mkYgCYTpLPW4TEMLjhAH/Qu
+0bpHz4jKWOq90kgOgyuDJv/IwJukFqSr8jzL3j/xnCDY86lWP36ovpByZnfJGoHdl1K5dni6pZE
TPRikRCywCdjyaF93mVTfK6IWY89C1QZmgMj13Mc2T0U8pYi4SN1Ebe05MFXZ/9vQcf3UY/KbKgU
RS/tKZaCewphAFJKoBIlk0YgOlC33YM99OtKT/DKtFDrGY4zyUVWYJY6C1saTmsJxQio6NI+5kjF
g9ObbMg/dtpoCaWtMFtvfZVQo9F/XWPNoALx+rd/yFjJmg+PgSVWnUqVfVII+4Jmv7F8fPz5rAg9
zUKuFgzXa+B3OWG3mbSIeEk1aXm4EUJorieNR3vZEOI8D0PeAPjnqIP8xFaiNEEg9SVykfnJjdfw
/tsbg07OZaK6qbSEqWmkr772+u1sNTEoUoIQX1gofAWMg71ziRJjh1IXFOKImCluUE+l6zBWCt68
vEy2SLOny0p8vwnn1cnNqqXKIdJEVSXZU3mbjTIDGjsTJUGtceR/IOLfGjiD6AbUScNH7oae8zs2
G3uye3HhknQ30gXaLptSehqNnpqCu+0l4iaACb+f0/CF0rB+ddrNdM123h7jkJOtnF5WMt2mfn/H
n0Uv5OQ+EofQYokbiX3brN+2V2PL+TkLKafmUrM+lgda6HlhVS1YEEAnWkqsLvYsTUH8/2/rpi8+
/Nr1z18UoCDogqsTieHkcSTWcbE8njdRVP26rGQ9j8zRgx+HOdUR9sisVOrL6yj6ZQQCLwnPLs5e
WoHNwPLW09jD5qFdrxtF2d/zJbUo6cMT4h+VLuddatsp4P0w2hsYyyQYxJb23L65Lea2haYObtUw
CRZalvdes/R07T8nLbTxg6WYCU2UUDV7CFH95pqYG0bf4OP5KleN1VFxkmLVBkjlxAhrkaI/IwrX
7ioh6QuXuK6M17/l15aoQbk0mdeMB+etACt7bSorIg2+NHk9Irie03cC1eho5W9qRDn2O4XYl6tg
Fj79ZYM1DDQ3qbUVpCtA5rhK2LH5lrzR82oPag49cW/BgR59W3CwaHqfbLBMZWDYQGn7Z2B4NDkV
7+x2SrdnYVi66ULacfH/En9q7lLkmXLNAtGGooh7deKTbWzPbEi2P2oqxb1YYAwIQjGyt228Eh/1
RpzbkrQYx23y43WytdrDXrW9gqmsfOB3hTg++DEYyJo9wkOjSAQ4JtgNLgo/CMbOgAC1MB+eKKPj
APOvmANfP8HhJwg6S+ZQtQM77b4I5VFAbOa1pMwIz7r6DcKiAKCAwR+bUX56xfGiysJikmIZ7LLk
WczCYqOxbmrfK2kKswY4Wj3Bi3wjaQjNk0DoYrPTYW+nL3GyIQBP4Gpa5f7iJ7BTdmGCDuL6WDcF
v+p2Vnz6stGXrRmEJau1bOPJFte4t5xC9q/Oohzf2fZxfYOgCMzwnP/GGhpaA5ymZOdmKQwE5c9H
MxtOQbL20qCrAXWSWmNosuU8b6ge+Uvu92PaO/ONkZ1fQLedEuF7L48UH/5gFSea7T1WgGtrkDSe
YXEvTgzH89zHQmlnzfhZf4+rRWq19kfAJQHiz2mA8xkq+AqYskn5a6049rpmh2i/OFLF6e+4V1Ct
ozb8bbolN/89ueEEW2aMmPmyJrXltkh78sD4h/Rub/RfPriW3cQXM5xIbEKkr+sziLUM7pgGuuJB
ZD0c135jRnq6xrYfeIDIrCWqRqrDrDBVPBQR9rAqHGirzBKptIKb8ce7bCp4iXV0PZmrlGsu3pSO
NaUfiaRdaRsWHQe3FXSDwECwNJ3zvzUNT43pUZFy4si/oXdPG82Wxef+5M3gVFqqrv9vasahDmms
Ity5Juyc+5JY6M1aCCqW5muLpIU5o1AJYpnba01LnkwJSh/m7Gsdluiz8idAVn2e0tJiWhC0y1zE
+AjpZDzzrrNaNdwLt4qdMZiEYnQ+T2RwkNcum0Lo7H/e3Dz63SwqkezS3pgavPK1Jh8fkzicF+Rx
99wQjAAOBRbOJh0fXWUzKgK9Dt90hwjMBLx0fcMD2i3OI0Bpgde6L39Jiz1iZnBYzMwZK5nhIpfr
Gmxdc7Ln5/j2yoPFupEpmZjHTLAOGkw1gzbAVdaMuloCZKfcFhZh2axCSXhXgNoIJ53DmFrWTi+X
4b0AtfsXxctecBU6n6Oay3WHuOMen3Y9HOta3DIIp68dZnFgofazaWsK6NuNCsEzRj5XMZkqBKZg
vLgXdxjn97+08Wifi1MXiIlg5G2F81EQgtZXly91/CWuR6iWcTCFsf1B46DVn2c4wqU0G4ARyRIe
1jEv3yBgFiMVzhlZkPgy2Jyame0u8EN0KLo9gdyku6/Gnez43IX4lfr1v1pLT229mtbF29n3iDgR
Rc1vyKisW7qY8hMhvmgEb4G/BPJhpmK+xEAMxO5TIgvKgIgs5i3g8h1DM45pkKeihNrrcfGSpOIq
AA6BZSPPz6VYetz12gs1FqhLYYu6Tpvmfr9qhSslkD87dx3mL2Ijo88UqFzWo0sfsxyTq0mAN5M+
hK/LJxYgZ/JBbzKirucQM/DtRlYGGqn2qJ7y9ozTWpdcQSW2wNcXQLU/ND0atnOyaGAavxqs/IwC
VgGBkZOeaRWtl0VR+NPmBtkLeqXbkSS0Bbm9ofDwg4kZzvVm7IPdZZd+8lYICxCCr+V19X0lqhHz
ezRw3T59FcPo9zr11LUdJd3f8577aABSXgVZ1m5aqKDctN2iRknUSpIKJVIuJwD6xRKODe6EJiwf
boORzun+yDsO4UNF9mIJLTR39A6jO+eZFKHn1gNA0QJVLfoFn8B7gYnGw/P568HZ+FdvL+hgov12
K1avS+IvLESleIKM486rtejw7gQNvpwkgt71T2duC3/n2TKTpaYbP+ToZ0gLkKS4Fa9xVCJ7NE0V
VvoHQ61TqDWtEVRAHjBUzzl0kFYRhbMOYk0/m7zBRlQNQKNL/BeKcxUsmmYlcO6U22MFFzY6qC5I
hNa5yUQSdN9/i6sym0cnbM+g3DOToFAc2wsjQCn/n1uL5/iTxUx7ycCshGfY2zIM7cwxZ/JUM06/
3vBVXkm4JBB8OIkJ4gN4tXvrh8T++DeOvdeM35P7ZmrAiPnY6L4ZOw2yH7r2aA9OSPDp02QxtxJZ
5QuQSpyigRHvQ8gvQSIHA7t5BeA0H7bh164oU0VERAvzDSCWGSIbkshMA4TgWnO67ehEAQm5BMIo
OCt53C/rZa4tST0klQKzeasJVg3JqVsioaFDD5A+sCZycRPgsjF4Je9VutKKkL+lFL0RXHcv9eTS
EXCdU2Q7Rg8hbGFR7R9OU63lDRgywctczt24Fjax2gsxHIRqHoW2uZggHiX7X0zY1VLvfLGMb5rQ
XtqpaXQ/uhggHOZXnIcglXjuiiXOEGRfkfQKqGLV12KjwhC1vOG5zwTxMEXKUNpOw+3ThCdnO4vo
dSZhoduXeUZchDGb/ciw/gDbGqlISSvTK7kzGvrsoYWRwvccOkwroprlo7sfjVg05Bp7DnhlFU/1
+NN16yGOvzwe/R+/nM68MfKrzLAaW+8F/OKUGC4C6gMhDE65KTFBz+mBadBxMi90EDTbe66sg7LI
Mj4uGnRkPGsjtbHvExDfBmvjwcaeHHNYmpWVD2opp76BeSp/QkbQqEtLLayJGMwqUt5VCF+54b9e
hPjdSZR0vXY4S2w7VOC6nO3GCbkomsfCEPLDvROX1z9mrfS1Aw5upn7BpTEI5kavNuGWvs38/8E6
PB+NWBHGRAXgLyKmdXNDBs4kzbBSyNHNTxbXDePb7/nEozDeehhiMqPysLU4iYOepEo9fjN8PGkl
OchleEidAikH+6XOtaqwNN9tRiR7/SS2lcRtXcNqWM+F8B4WVQ9qIg2341wYGplW9/EHaBTHo1hz
yWYp+oJMH9Q3Hl7cQ+jZGr1jKhDv1t7RIOoBS/O8KQ+eHl6YQSLF06vblfDM2+OHxjRL1wVA0nPN
p3kmrHWRjYqwwAbDHqaLuwBAwYZ3KxFDQ7pTWbseoufQA52AGdTtHzIUmrnNu/1yqtr3w7MQFy+y
S39ZY/9egbHUv8h0scqraygHFqn9e+Ar4o97pDBtxFsnBDeEwGBcQ1jd5VIdSVWZXBoZ/Lhp62OC
iRNfr6T86mcCcyTRhInqsMW1tUnWtVuQfRJeMBskzNaIWvwOuJogxuosfn1kOGeCjTqfmHsy2/ij
MH5Z8pRzZwyoUSpO3ItRLr2Z1R/RdaLRwLsMjg/MlsnjIAriOnoosHX94lJ0r7OtTgAJMdBeLKCP
a8X4ZJLry9GzL2shQxyTtHZA8r6T8QCohgBfF8xOWBbt7H6DvfOj1RntbC/+YE5lEUyXQZeiN41y
+sd/DcWeVwKz+/xjniam6Igv93Lz+psVlkv5b7A5BAq1/XRpp9eEVqY0JAIw0T9BEHTUGy5WMXT8
RoHwhjrPwieiQmMjnxD05u3uYjYBji2oWrfi6RQxMG4SuoGyWpTZnWe83n8mkahcEZpzkRA/AP1a
ubu1HmMonZPVNUD2TfqhvqlQ+7klO0z6RvpH/mAO3GjsUEVwg0b+pGnQlwnrtq3HePb8JrtnfVHf
DcjtzE/O8uRQAdFLLO8tqx+8s7jBFgrO0hPURoqVl1l4R2AwM9lKKpmGml1ASVK6nX3/CTmCJM2j
OMeXX7c4FXKSkuXrXQYqABEwXdQLdKbNvEzVe4gpLZ05P+ayNAy7rZKV5a9tz8vOTtLSUvSrLAxU
4neIdOthiNNXO5eDAo1dwFkJe5pd2f50b2bBlEn2LaE0aoQCtgF/WIpBIQuelFIhJL08PRzkPQbz
tawfftba6UHsrwaHPIZiqqsvFl7DafGlvFaID64MatL8iUzwoTonnWg/neAoeKG6xG//+fpRysN6
RY5YnBZOz2dXmERiUjE9qley97ikowJLENLhjNgnaug6Amge2T7uifjx7oOph2WkEuoWXbsOE5dq
c4f6Ku4ZnQQBUmBkkCO2ctxFjS6WoSCobwE3qngAuGHZ5msatyo1mWy06gtBdVXcIcPNQcwJFb4x
qPtAnDoe/LANFL6PPGRYht121pWsbvAD1+6LdgUyUS88SQLdUfOEByfL1HnUI5WCb9oE90QXNBs3
gkvZO7CWTLLkNr8F8NvlENZ5fAO3xWRSalx/6lONFN1y9kTcERkbK6XsYJnC9qT63sTOPABplC4h
+UMCvqW3oLu0Qzsrbn+3LZKOWXGQ2FT7hNqJxCWHc896LJYhnFruhvSQAucoCBGPqj++3AzXopgQ
fOxddj8sMulLPAkgJ+7tLEk7Pp2YW0bjoZFdZjnETwR1jkUvVgWUuSiUsu3Wb17fjRwdm0zGwrLM
tcBb7J1epPUr5Bze3s5bjwEjUpRKyR7KsoYkV+5FgoRlvQqdhQVp/NRVp7EnA0RfX6pDEM5WImLA
PmTuXuKezmgRniepyvZeEC5T+JRonIfV6SLuO/H48TVEt8eJRjStF0OVmwuzm9mAZXntNqfstw+/
klj7SjnmOojM4vS6lrFL9DSfmQFE83bBnyn+EJ0F87zUWCQk/FiIgnpZFx2toKNXjEVgtx2Fkm7X
FIxXUppXgXJiZk2PERML555pgKbmT00LxopAZB4By1P1o29cAmIhtMlhLrgmrDLPct7158aQEyNK
iRK4dBcex7Jy/IguQ1u+u9K1QS95NWhldD+c4Ng9kXw+rWDFndEGyBaS/epcySlNHgBSYM8eTRpF
J0B7nID8qN/M27sXfFSSuB+ePdBoGrNhFdVPZLUQiGrikygnzcgpmm/1J+zj147dM+cjGsnb+n5C
H1G6JI1Yc3uqXEVP7TVG5GxsleH9a4oMqyytPrMBg/LxhkSAj83wr1w3eZo005y8RLrcATeMEDTc
8xR50NCjLnKJkARhfT9uLA2Q1N0nwB1jQsF79XghwaldGtvKK8ulN5f8Hb2MjRL3eWDCt1XBgOlg
4rbgWWqXx1eahmNErcR+B/6GP0ErTWezrA0XUrjgmgoF7Jko5KH0Vmzw7J+zH/dBiXhppUNb6Gmm
zV/ubmTXYigJ6HZDOZMxNOfRwapGmlSKG9gfboqPtJaM2yNBw5iB/d83u9sJWzkLIBTQ0JMmkcUk
5mrkBPQZ3fLyflUL+JKMPU6P6bP9spVwKecfSYtSeS1oDmuRPogP0CgUnl+CvR2zaJmJbKadm1z6
tBqjwRzIFmc4Oqbc5Eb+O5MUiCOkGX953x+5YOmLBTmQoEQP0zKQw5soJcv9k6m6ilQNBbxu+i02
lOMRzgAWJxcKg7PlKz1KmX2qatPzt8CBj0XuyBG5Ct3RMk7ew3J3LEWUJXBp9aU7rvvYK7ORxYIh
4QdDK1od4W6WKqx97hnwau/tUTxSlXvGt/rseeq5B1aQA7V09AKufBDO6VYZFxeItcbuOiQt2j0s
3dWq5P1DFSy2BUYJPegTfnBqgBniZ4ocIdR53JUkbtcz55mE5d7g8y2boylQ6bkpMeu4xByyBlIM
d0DoMivicEXw8MMEcjhENrTElFgfhpvB46jyvRk7dZbvf8zVH1H+npTuxafl1zgPZAOLM/8IB7Bd
ZhkYyvPTmJ+9wUuLlYLgKNvHXj9PASfENXoNv/E5ycKJCinsuQGyfYTcNcFpz73Wolg6AWNK6rlj
dIoSOanZ7QKMxyu71S46gYAWQGkuaOJK5Qk6lYYrRzqs2MINadDTuTltLh2CIZnWTnWo2+EmE7Zi
jMvqd23FKW05kUNEOtwZdGgSPDt4eBqT+4xptNs0p7FLPwwMQVD1gUgo6q4nIXAsralzYAFzHfII
As/wlVVrbxH4KejJCN+VbOFs8RUYgobHMaej92P23qmSZ9cVn6ricflSP+tpFkdQSIg4j0notAzE
nAbITT2rpmoD7yQqJSSBQAyXaMWV2VKsNXnEIHNK4db4PInbm+USA44XetPDqR9BIZUQPmZEfmD8
s4ANwmowvt99tl1lZ3g+1xA03KKcMzjeUSyfRGL4KWTV6ELmeNolT3Jv+Rr3TjQO8tY6qKBqJUH3
7ZMOdNo7n39MZMg4dhu6nzlpa1zsWugV1PwxtA8VLQTk2MrfH0HgqWb764ERWIRbWS3KpDXwRXwg
9T/8Y1t4NSXTJ15n/yyCUFVdNpETWpxtm7F/wDnZbx0s8M4SIHr5zT1aADRHir2jfKHw0tJgp5TG
DddJReLEe8oBgedsiBoJ6sJIy0/4BDDbhxrpOSe9wzGmUjihafvSeIuT7UsVDAs5q8FFjxvsZqSX
+HMUT37J2JitoS9kWB2Gk/HT1QjDyf8UbnPMu+puMgQtT6idha5lLDbn+mPfNDwwVc2SqSkAvPjb
GpMv1F00TY8r19aU/VUSYe5+oaYwro5jIRXsIdIBG9ovRBfJP/ei/+T1HamKbeYaALP9xaiNFr4I
6kxvSUWof5/p1bYgQYBfIrGAlXcqdTa6XIy8Ht7/rr4ZjrfV1I6t+S1tvrtJRP5S1lNH9oad+RKa
aCSXrD7pnOUp1ZdKPSDpBjdwE1R6beLlVB5XODvlcBS4LDtuyzRrJ4ETeO3q36CkdveLoM76ejDc
QaPiC1mlHX0OguZgvr5FEWrjJrmxJDxW8+ZoZH8qiw6gEhWvsQ/TXjOcKT5qqcpac3t613sBvQ6I
GTVmA5s9dZeVK6d7lX1CquX66i6VA211aZ+B7l+TNQWr6C27OljsaygnVqImWMDy07tL7EXLXhSr
Y7BV1Zg81vIhiu1jlXsCnm6r+d36iv1gJfMujf2uTCiq4PZ5gYPoifb0g1muIgbOA43iRtHLvHKg
uWdqWYzit05XZAXyYVT7SsjXvmdiLr6RjVcz1Ens5StuEUFMaxkk6xjR7030/N1AdeWRY5y2or42
AfEp1FBPI9jJiWRwVjLSP8CKyHNIbv5jkqzdNmqERKijlTIh9bzqF85WnV0MTfhC1A9sDMV9sTu7
78rgBLq4yRIc8Bin43+60Tawq887OMe29CU91R0sVEUmZuEYJ3rTis4a5TMCJ24XeWcc4VGuyJUt
uWdl5h4i/t5T9ui4waPrn6Pd8qKDBZ3U/Z6WEtx+kXGeLTXUIZMV12IUFD2K54hXXTtfFBbhxnWZ
Gm25gDU2slrDhdCwK0bgr4JWr1/PLT76ggzR1dUpbfpzR1E0YW1vrQ1LTFqX1yWJQv7gne+VaMdM
ftG2fCdRUEYm71QpR7qNQ9jAlVIB2n5y8Mnec9kD+0+dOiTuZtnE6HHfHnHHO9SMsmvHZy9t2WK+
IRXK6Seou+D8tx2AMhSxLUf//p7Q5s+hbzNbjrrgt+bJ5OyLbajPc4DLplTnhXy/IDpV2I0kRcmt
ARBYy1+iY7kLIHOPDXmSLTy0TF/0JuJIDAc77oIcwzhefKPh7P9QIt56ym7zvNftX+ycVlIj5x9f
LSyH+fPy6m49Xcnd36O4rzi5oJ9qgjL+w96BWs+H9cqp5goaDrQ0o1WBFHIhDCwFIrv41lKJSezn
c9/zH+a7iwq4ZRZ9BNRONiwP+LianUgqsH5rVtTUKTUiaJZocDgoUWnYSm7Hgucd+4JXTdLx1wWZ
M8UnY7bN/GcYUBMLHOYD9hBzjdLE3GjbdPP6Jen3qYXdmU8xPEIjblreBWbcBOBvq0bqcLJCA+wd
8y6Zwzx8zeUNR55JTPutPUYuOlj/2s5YYBaW+a0LalBHC+6kcFdgGLRc3EqrbdW4QPGOTdLGpju6
IHpkwXPRwzH3VBXwMRaYMvEkzzArfGqOU9TEIikdXPe+9pbWB6W1VQoPaALE4QlPU517Ru8Ia7uT
oN0CHs/iyrjOlicWnAeZ0PYKc1vNyOGqi/NFeI1uWqEh3oU864bFJMdeA4wCcwT6ydnbbqhftCEW
vmwntp8F3Qhs3nwhrH+iiwfi/+/ztXbPFDMCDg+nRVjv4Xitp8qUKJnK+gjm6lRQt6BPr+heGCO0
qpwzxNc34YaZPXZoCH/xDRuqNcWtwbr+fkeVIbU59FSVF9S45RWlJEOSoa5XO06x0Cvu/jsG9Uex
xP2FmJ9xMHCIrklk0XNN+RfyQOp4IrA8xjMNl8TH8orY+mjcdC/26EXulsZ+bEGKRjzgGnlP/lY/
A0xSiFW2Fbz7ppo22UceD/3CY5B3JNTndHhdaBH0dF6qgVDtpgY7ootCKXZaLCzSKYd7rZA/P9St
g+vf1rvKb7sTv4R9VpAXw2J5PZFdXxjk32ZvnP/WW4N+hzwHGRYheiUzuCdjNGhPpANqXuaHaylD
Dpi9hXEU+HntQCHWMq9uYo4D+yJtbqR37Tv+ItwHnGshRizNMqr1fszso7Qyw9iTkAIH39Me5P8+
tDaySOqTFRFO61dS+2mIhZmN9qYYBMoZb3kTCfdO99eehqHbYhnMwkearwZAmSLlszBD3rsfUSsd
+daoCbx0Kj+uQg2YWZJOZlIg1FZqobs6QB25wFkU+HzebjrfzvyW9pS8a05E7ZXjD+HaghyLW54i
bH6RRZIpqzZ31rR1ogRjmf7wSQgVlKz8J147RQFWz66mH2UNwEK/fqBxDdixdGZBzD673GN5+hlb
Ux25z1/wCXv9eawiv1lJcitsf8fEJoCrr6zoJbt1rZ5ic6G6pvpXh3TC233qk9dNHFrh/3pSa1Rj
Ss8MsILV5IaxCQRFOx7owdo/vg1tNvPaXtMbHkVRkqc/6MoiF86A0w5PdcBo3dltqVLmxhnOaoDo
svFTYsMahOVPHp4tHLTziiynHarDiQrRSnsaJ9tJjw1IkbyQ/01Sn6gRG+BjdjVsIJbTol6oNb1o
M+575oyXhstZz3vlHg/8eqd5WiNOdUZECATqNN6V8YV/l3woToOWrTx7DHHfmUtzwcpHsOHZdhvR
EyG0tNPwDfNf8Rbsh8hytq1plaQCvfLdvQMTLwVDL+samrO1WHdtJjZloC4Km3iuNoGm2rSdYiyy
Pk8BtsqEI5meSDg870jCrhmpn9eZZ1EKcXfyfgLmNZggHuaosytjC2jrrQb5O04FuydSYN82ysjQ
Q2KjZ19vM+6Wleo79AxDs1ygkB8pmQ5mpV/ud268B6BHIkcF072fTj+YE5XejLV7IjD47B5KiSLZ
sgEqm1kuNYXGFxJCg+jAd7d/7zJRRi42kMzG2rupus/4b+Kf26mVAbGKx+Y6jDe0abRHWLTknMRe
rEVNxZ1/9X2oQayQ+UOQLamfmZEjjYpdQOuGWJ7f8WMM1nc+FyXy43BRcn03OnDA2/xSivsMenud
kwCZfHaaoKGjGuRr1XkiIxpKTvkoY4xbP98nX050Lv6aHhiKvPOclQ6N6vTf9Vl7NZ+bF2RaZasp
V+00b0syLiySfp5IAscL4Q/z4SVUeSOwXOd/QVu75F4w/BzVnaePZt6SQmNv04ISbB3uBreLy+PQ
v3Oka2yxUvVfxZjZjE5LA1dymOXU9ZU5g6zyQJFCVCE6EVYf3HbKklUVeQJS59JzMjBJBxXxKxdo
FaTZ5gYV2LUWakHEvlN4vsHHslPsuJpwjg4X9MOg+/YwcpFPdx2QYfdWsMoyiM5v93TJQ4EwM2cX
KsccN7HCd/RWM6cGjgLMBnlWGq7GWZqQAdcakU2Phnkp+KlrmgqNhWgdGUcQbnaJVZNefl7HNcmx
b2vOkT61qQcVzwyGZ2krFvZEhdlPWVJGFegZ1NPDwyT086+rjzlXx7t4FnDLcXJfVpHwBps2tN6w
TCJFXhpDtSWaDhg/2yfnK0EklRKK2a8AFW8m5ZLQk3BsVLCGLNXxurcusxPUt3mVnzB6DyY0/M6C
26a4eqaE/g8nsQcE/VBQboNRicSCX58r/hA4kHRla9nkYWgOGDA93aYaj0dwjMjw4mruFelY1V7S
BAfJUfqvG16Xc7/UKPhRaSZ+z++GzkgpCiPG5ajR0BdjGnpBvPGtQFlbndWAVpCRXVTPfnEfmQgm
mm5B6dtydedW6yqnDXYH2Fo+/qXYLS1s/9D76VUG7SPoAmO4W4kqCpCSVwBqRBHK+TRdxVtnC+hv
WaWr+yG75hgbHafk+ayMCB6dUHVI/uLnDX9c7oJcgm9N1k8yASz6VT8s8FNckzjVrcD4k7Eu5Wbi
FsIgWegzhyptb+rlOFp0yF9YVINBg3f2GyXNVG9Ceu9OvaJr1N550ab652oqaMSHvpvdz3QnbzTY
btr0MwCNrXfFz6bIJk/ugiUCzdMrRDdJft8JhXn3zKQRO7K5EiPnEfSzD5TFa6YlxsHPliy4jG/d
wwhwuL4RvbJJGLqCVw1oZXRsOhVjet4gcc7xQGcnrE15RbBCitb+EODq7HVggY0j4NuBtwq5Tie5
OOuMSWzdesvHgutb/EEUlqgXpIEL+ilrQ7dibU3NGEJafVfSiPanNz8vCuFVBhGRjrdmgSNYkQ8h
8H+21fGfZYkSh3wVNOkQx6XPPz5VN17CZQi9+IZm9Tcbd0z6SHWSVHv6t6eQAmCwJ5WowEWmuddt
DTxV0HfdQ5rJ6pkTa0jX3qlZikwMk/f1VQO5vi4L+++96Cjs31PjG8R/T7mKiNOju9hf29aKnLt5
d05eOtahy0GK9XkB5+/+6MTpZhhLt9jdgGx+tVLrnM0NwalMuQ8nuqQ7DCwPnvsxjbXsGqWRno2i
w/SuZ2zsPZr9ZEg2lu7ywCilKy3hBFmhh9Ioik6BQMcTKzVEiRs0zU6NM/cEuvh3qq/ckfKsIz2H
Y5DFn7ZdyDiFeTe9/uVs1ZcDn2+xCsPBlhdWM5MU/0l/c2zmYGazWDwmFxoWtN+qr16b4TW5be2W
cmKh846rDTmbK0N4VaveNJ7hPaVfE8lLOrsenvNfBDhiPRyLvJs18M05rLBgiGq95j/YiMjczRKn
vxRJu8Tno4i1my0PRTVWBSX/mJ6eacJYyvGnJ44pODUJ0vqkC7gq20HcZrWTN2oJbiOw+FBThgbd
fTgwqRP2mEcF7rUEUiUvbZ9c7RxjEQnv3f8mFxdvGifULNA56GQj8Rv4UzR1Ha/2IMPF7V8qVIRN
bOuUwJFwdWthWNl6x3CuS73pl48VuaUnKMEIHCHThlsWDuL1YJpH/4UDKMqGl/JeqjtfVDdKKm2V
jvi+m2xSoWZZH2GPL5iqGIXtAs8X7oBIPZuLKBVXemo/LP52L7TIeSmDyR41KfZpMroZ7TPzB6X5
DIDHmza7K093nSbbYLOg3vyKFQfkEr9OiesJh1QNvSEx8OuBmUhqCyIrQWdOdNk7pEHvEaZjvyD7
L6pUF6Nu3d8FSSOya0hVISIn1Fen9173ne7kGSDNbAJ99ZXfk4bTe243Chv7+Uei5S2batXRnA48
VGU7I+7BjkqAiW47b1P9lkmSAc8nltdPGx9z1zyPwgKET3HxoQiL03631OKrvyvzg/7kod3hHdNu
S+sLDx7Y35GSFLyK5d+SACvXPqyD1EqICA8XUidjkz03twTiMWEdRjqpEYMGgMxCtqr/qUmliS4H
CtQPk77Lkl9roHWb302RLqtp70uAFToI8AB0E2ZF9PzIWzNVKuLTq/cZJGBRp6vZIYAxXXwKoQlq
B6rdgJBVOE6hmOK0/qbmjkmlndn3xQtQ1ASo6UB+9qabeKwapi9/rc0G3qpfArPxle/qjYdRTgvM
biSv9gLe3JtSTQ2F/AG3xsRD5ejt95gGPHuL4B/EtKymsKIhdaG9W0mWR3myZpJxnSjzWNm5TzDG
gwSqfuFIrqU9Eii8G4SZt+Y++3HMlvpR8seUPga8E0aL7Em+FDGccHf6a27AOAm9Jn4uCSbLiELK
NC2Qp2s7xfaQtFWPLGqDvE1RUKr/LiSawF9YfTaFytiTuuOc25VIoGvMmCz1hQc9FCjCXgzwM50w
dDIZhhE0aYuSxG7Fguoz4lFrs7IQEGd8+7UlkN4HI1VixIG2tJawtxtNTOfniIdJ/AmA+aexSc7S
5cUkezHLzoEPS4DctNEcOYGxzPGSEFqncp58kQ2/Q0dRUFJGzlKvxp6avNcWA8FhV9v+A7QNg3KV
mIi331Hz/zEyVw4f4gHVRwjsd3UfJWDs2uGHNhAyLJmACGL9jAxGxSdaZDPKs8/rV55lREhuvx5b
BAP3ktoW2BYJjHy17W4ik9bPYk8OF5G23Cj86SeTTMkQVG6E2AXLroHX4ty+o29kkbycH8Xov7lK
CpnioLpYaH/ZbPwe15MTQmy6lsUA3VfbEhPZFKdhbL0/XEG9SN94UpOs2ufa9j+RJMR7SL8P4mC3
77o8uBv41aSzw2WCyRlLsjuziTKQBjMeoIgndBDsKZvAWLXrEGn8KOFFqvqXvR+i1uSWWA1+ueNi
38yvvEn0n27pbT7pMlQRH0V4DuBdDiQLQ56iwMMfr0kWojH7j5OSsrgKiwjlSN4TmdbbdzAYLY9C
mfORbcSx9HPzxctk06cloF+Oieu1ZyU09/ODzMPjWVvqH7GVDdvvsZmf5SgeWWdPpDTRNhPmTjwL
v+kUPNjhj3quDQGSpUWuZif6wC5As9pgBZNaATxP+IwX+BYJi68fUR4QHx2y6kXogLJgt/4B0QOv
SVv+X6ShPDKwXvlj511guRvIR/fdpQwSPTmpQqeL2t9JfYhGnPQ4BEpAnzNVDysZBIBZOVUIiIhr
pXp1fFY4OYGmNvrom2DkVNcUF4dMkkLCD8t7sGqVhoS1UO8b/Rbhw8sL8SLLXSTZd6NKK/Imnskp
HwSubbrWO+pUD5oztkRkjQILAsjjJwcEVoBGq1Sz4BXei1urk+4R0xYvAeSa/JgKN48jVGMspcB0
Z6o/o36L4IrIByxzNOaGpBXYW6au74b3AdZgH2CDwOafN/Rp2qMabmuYmkm9A52ZNkMc03sxiFhE
DxCKGmqMsZHRocHYmW+0NzM+Pf20CTdV7REx13mva7auhx42DqRe1TVaeQq2pH96G3ikt0Y2yrOp
S3Wj9mZPUTQolVF+E4D9jeFYAEI4Fsxw/VEvEi55C4zyvkOBK/6xHqo8plSN8I4zktwX1V2RCKj5
UITUxMDWN97CY+iZpZHNjQBuC1ftk+hS/qsg8K0JmT61HTUKhCBnXzZO43dnw7u+6amMb342OYtI
IxXxsU2+lw0huR33+qehUfdZTf4vM8hDoe5IvydlyIFLw9wzmnmnvuS17kotJYayxsVIewzJvsaq
c0hkCT2DYDgbWWNC0AOhm0L+LhTmGSMIhd18t/1F8OhZkEpeGuqNqqhMXntZfpeR4wzGQNLp7hov
oMtIlHoD70r9NpYDcYwUkn/mxKvgKGGsUY5gSzgX+v7Hkt9VGUM2Wh3ZcZ9QWBzgNO7KRirMBn/d
G35/3mAnoduOG9bSc3BthkwndlKTbVl1yamw/dTkrVgAn3aKhWIorLA/P0uBj2p1vzivOAJLYaqg
lPHR8oC+mZcy3NLfK3CZRR6NdtyA5kHevgvBJn4mv4yO9e1ok7oEDX9+InHS9kNQgat1zM62gZP6
hH8xEwp2lns3jsDsAisDqF5P6jBww6pUT17GVT6lfXIYLo9SKOn15H4232TqCsxzfANI/dHb9AU4
iTzMWnkU6/kpOc3x186ZREO92jWd3R0n0xiuceLaPQGYZE1L4giLBbrIpRYXyNihF+A5Fprk4mYm
ais46aspxvHQGgUkX7DZUdxF2XrUqU+LsGIXBmW/F48Ruv5/g3fEumXS+8vQqo/XDTNHjiNJBpyF
1MULgaXHA8hBX05FV9Q58/9DGc/K/nvKjNLd0uLgiDLish4cF/sqNiA0t3kAFL7xrkoIUuBTWTH6
pxXcC2NBYCpiApv0G6kVAIWC+VSYYaaTM+XqTSF8r2y+OzvfLnXH9wDx5lr1bOaHuaxi/kaYzjWk
sLUgxUMjrxDPmb7yQTFdhSFESA4r86LaXIPpSkb778wC5kQxlbp0al/iiW4R4hu3sG6x0Z1YAoo/
swH9qASOb9BakBXfyl6M/xgNOhI9MfePWh7fRv/TEY/EcIUjfM51xNHyjF8/Ku2lbVd6F2OSNpYz
QERGDIQOvIyJs8oINfaPJrhiDt43vXuneT3uysJNrK5p+EQ5DxjHL25K0qH7NS7nuisejpW1PKwu
a2sFEx3q+o7a7bGfRN6BO8YH/Qij4WT7xW5CUVuDd5JuvMGo2nfpRR3SxZTWwfAJJUm5ZN6r2It2
p/d4GG3+TMTmAO3QoQyHGPcNSt2c5TcxMEpRF4oV3BgopZBgujDXsVC0QWQJJxRtfoZ0Llm7LPjU
Gjg2OS7iSaqipmlCRd+wh/RPFsMMR5YkqWMpIbX7koC8vckUEVoifrf851zQ2vMICJ0xcOcEFru9
zHQEmR7c+LVdFfdBQhujygiRIS54GEhiLlOJpoM59goKzcLdUCvPM0Y77t+Rw1azsJopxUS1oYTL
CBnd30dv1+WN0hr6huU4vB7hS2pz4OUncU+r2+A4krd78QeXyHzoUY1qs8mLVYEWmZ/NRdjDzJoY
c4gEt/VadM82NaAHdS6eEyOXfDWQzaC8nsm90CNsso8VcS4DwkIW5XBXIyADsOJPatZbAJ/y7XiJ
9b2aX7Ff8sHhnTQgD2UVD//+euXxde2QVprCFh3Pv2HeGrgnPPFihlJoX59Y0bBVZ5+lnlvKyulE
8FCSlDw1hwCYwebqz4zVxW8qKwxrYHrGqetUWpbPvI/B/NicexQqVsFv5kUu85W+iB8Z35Kr2Cm1
94Pi26mzTSIzkxWysAvo4nWlas6MbJi9HTT/Xb2M0Ad6L3TVv3mQNbkiBBwWNLv64I3ysAZVx7uF
hz1q/MW84yJKXnUQruKhW38XVYpO2ttlPVI/5atffVg+4xRUxbnyrzJP0N9CbU0ogspf+pUzsRRq
RLLKij7xfjuPa/A0i4KxbrB5TmbswelN1NUFMwG5bPzHw7jaNfJJxF3Dmib4N6susle2+4xPrH/n
fCpzTUZLCMqH74TvBhVp5euG9aLzjIzjzX/CWODX9xyXaaprL4HahZMH3FMi9aanJl3G7eRXdqrY
06ZsNAmpHCPiY6nvec5bBEZ9v/BIM+5AS6uXLv00lYHYNNfg8Nc2XXGHuLHkVXO/CMhqVcUvr+la
mJZVDczYTsBF2N8QyuA0CBIx4pY8UyZ/UW55RY4sxNGmw+JsEiqohrFk9zabaKftphcfOdC9FNa7
z6wSHd1pK1jQ+qnnYWUJle9/hCYWNDhyeEi6UPxWaZme3UlmLEuwY19aMRAXARdUz1wD3yjUCMww
k6hgnJk5dpyJ4LeM6TsYf/NrKNUeKOjJTrP1vXMuNB2ada778DeEqvrYojjeJgWkw3fO6EucQfru
n3E18zahOQi4IIXUj4OSHrRQhTJFpoRS92fqO0TpglxHL7SAA3mdiQBr2lqzQZnjknZ3xFW7mMTK
sBSkCM2xE4fhPsA+NGPLmdrOFZdFKIzghZTFInrzC6OMboTopAhruakiuAvPeGb8WBS0UfraaBOA
hMQB9znQvDlM71Q+r/ZEqEVhsA1dMzyidWa09hxmDWCdcxrZQouJJ9FIsihj5tTQnaOCL0h8/sKu
iE4yOwJ5YNueWAgSJCABHfi60CbT74IXqx2S5te2bhQcXPWWd6fIfGaJN3mj1Z+TsyiKgU48cPTt
iOPh3aFGMOEkU6ih8nQRpejZUFgNuzbRdBEqZaJ7juwKQCqyXtEFKibIuRnYmYNguryQi9IdBgkP
trLGbg+Eo7FxHylY+iWXy8oWQDhiKpB0fRrKLnpxfaquvX6dWWyIf9zB9FxVmMuueWlrabTgbtJm
IB8oUzj/MJPNQylHpNq95qKB8ji2cCIbhmgSdxfCKeax5AqNhM17qODs/nImQtA39Gw3usLMzyeD
UsI34qPodz42XFwU+AHRXXDqpbXWR36QStBK76WsoFQv4ygCOuIYDX1ri+OzBgtlHEDlRhKm0lFH
SV7SF3ISBcTKfH0gmQCuhlANqztWZwVjjC+KeZ2KO44FRI7x9x5k+7Co/TtAnKykfaTj6pYrXMSk
0EOypcMUJ7jxXU822/JNlsyyB7mxKmUDpJgZYvAFp+qUvRbIA55pRuXTOVJbGZRAS9N5JWGiArfx
R8p22V77+SHO5uDlEUO2NcnomPGt88cvTCxFYZpISU8+iNW5UaP/DvoAMEQKm8Fl3/H+oh5z1SAw
cQm0FRIQavUtj4gO1Yk7swCvCYEGlgrh1p0SanxCvL7yKL9S9oshWUqDpKvhiH5UgBmdzTCBgPco
lPHCu+NR1Za/KGBRgomHitfDr9NLxLtO8VueHf8cbVt+SpGMB6a6pEqnDhLfaUJGjHze+OJmJPiv
EzgdSi2ANGLQp56lk9C4UWJdhAYmVcYotYDLYSXj9ncYgMfV7d4x3pojyFUKhEgDqRlhbocpE107
DI0NVp+iGfpC5v7jgMbi6Bj1MCKXD45fjdFjVLOghbgNNlrXKQSeHYhVbLkv2EeEw5svZr0o+Swj
AP2tCD0Kxs1j8+BRGh2zf7eXFLEB3kFTwaWx15CRt9D9nh7cfc+oovxv4oovkxkJLudx99WNwxDT
formTBisn7sjTt2+k/ZYJZZEEhl4gGBwuG30n0KNpwqdt0Z2vMOqJuAVeG+oJALEKLpmHz8GcXDg
UhicvIUk/JgheMntMCvr0+dm7RR9KNuPnCv0A/2fmwWxb94Pipl9+5BJ/FXhDtFiRWh+6/YW7ols
IYTPoYWQyw11tJ+Jef3joG+TE1bgnZ/2LRjsQEw3C/i6+8aF5XA0xYFj5ZmZ49MTqRSe2gLaNX/E
KcdfEhj4GIKOusI4AMGdOKXvETMN96AC6hWHpceWFkfPdI5Cau836lkAjF8uKm1hFV5EU6brxsq6
oh4L9XFrhIS/ZoWyuYChdjHYEf92rvvcjc+M36bIwIyWJJ8TUz4NrmcRW9iNP0gExF2Tek6o1swK
ugfdD8rMnXSyNy8QSfo2O414YJG5lgGAaSUwRxfC8PYd2z1hP9k2KghF0n6rYGoVMxpwPrzR4vEB
/MEn5XDE8KxCbjuOJMxOpUz98wJo0CmtTP04TQpli1Kpz2R+D54NKy1UOxDt7YRX55SGel5nm5nD
3nPKA+bJPMW9PQOHidEUwdU7qm79EDCgMjQ6Z30g4yQfnlyr4k+9mZ1qPN9+Y6qiBU+IbWaCszMj
b/Rxjsg2YUXwCKCBGSw6boXuXyeWYV9ttz7OPoRWxGUSfs19UQ0wua245d/HO3dOHSOTSkgMSZDs
FhNsnExuZ4HA8rtsLsgTLXAUzkNMfmhQxakE5SLzcgWf0gjaETeaBflg0KLzKd5mHnY5Nrx3to9/
dMpYPYzMjmRIve/SLJF0rBqT3kGIHd7SWkruEhKpPmTf0jii0FMPat3JT2pJX+M2iLFChg0lkzz5
z3gmyJndkxawVORz8ekA2d3sXXBeZ9u6NbVfHCrO2hZnGnxq5S3AXBxh8ZyNz/UpbThe+8r2Q0Jk
GXqfyYYpiy07A5N9stpWTPUg1Ni0aeGl8XjlxWsLpBdUHXdkhDp5KofT7Z1toQOw4nKAbzYZgxv7
0MutixKH4iKLgA//cYMSf41/qZFVPe4j29b69aHiNAyN1At7gtMiLMWfXf8zTnyFJ50AQVAWVl9x
tH3DOxpn9F+voZ3xQLABUAmlp3B77DsPeu7WZtshWBbAwS+zgYqeJ4Tj7FAzwDmNJRaYEmAbtfhE
+OdU+IT6KIhNbe6/wdoqJDWIPryh1xOq8lMXr+61TEp53JnvFuZt2bdM5orm6Kn7sNtOoPJuDACd
jQ4kk/q8eSR7jwgRZ6WOwoi/m8+3+nxoRxpSIN+hQ2kC7F3UE5UDaWm9DccZgcmOrV/P+ePJcSyK
pqt/n7h4ste4G2u22kPmcR58qis6ut/duX9moxRq/qUG5if+ixqwd9DvEpuCtXpH1tsUl6U7QsNx
t4SAGwLI4UThO1ELyoMnzD+qttTHrroV4uEnfUpSmr4LXgYsWLjgpTN7Kb56PDTj602HloUouR0s
YQ49111c2NmjpKx9VDrPJIUgfnnJHm4f5JQ0mgb2x1jWq792Vl+b2b346iDM8/dg7XjPnVLJuQSW
MuHoPACtPYXQS5bSTHT9wPI1AEoKcQ3dId4qONj2Cg9WrjPiM2lRDIlRe0Zji7U1eYHSxSErObU0
y/Sp0cPo7o5rt7sMbVJmeZRajR8vcuMzJTzet9ccTsf+87UyUAYpP+HzE+G8k/xbyzoqy5jwQiNL
m/brN9aL9rKRXjNgvL+vwty9FuyfTtYnx0+Cbt53LCqiOKNHtruSwz6fJ1PSAooCf+gBzCjDWZL3
ZMJMIUgsS6NPhnQhZV70Mh+Z/w6AVWYeOxRvajnL5oVeOypw8tJ6pHz/pYRh/MjASbOsUCX2wgjI
PWDs9rCMNOzAvXiiPICL+6SoxpRmy/CxAL+9Qr/vNG1V0uPCfK6T6VY2RKi0iX7OcZTIZuux5Ry1
7HCXIcaxAYlVDVx6S70Hpll1RKAeq7WbOwIbbmey+GsjpIW/06iXGi1+cAlBezo9EPT7byJHtvPy
rR3YgMYQGs7w35zQrZT/d8kncVTmk13s3Xs/c0yBzuCiuZPRb2/oq4tl+Tdy7tsgF9VNH2OoqUBX
8MydaseOkkVKIuEuWhXtuyy5ULgHd6qucES23kF484GvEXmaA1ZxW2tSqgc74qKAlqT0jNnDIMtM
ns5a4bqd+k0aYEY3uLc67aMYnp+tvFm7SYypMhcMV7LEN+3x4gIp95fXp6RDgPSw3ER1gW8/tKEY
3Hl88+sfz0uCJs6rbrc8j0xrh3+Tb5JxptYQwfxG84tiSW86RQlxl75Xke7E1g2Ib605kK7gx1UR
ED8bJGLxi9ILtD67dstZIEMZYq3Z3Gn3bdip95VJJDKoVNnSz2nDWhC9h6gWb7+w60nB1cgx6MvG
8DyCXUAB5Jy4KvmXRHY9JMbObwV9ZePG8omDAfnchsKISDHv3dYF5/O8jpVZBQqSvpDQAfMmWcZ0
bynbI4g641eaKQ0ZkqszPmVglEFhT14rzczMb4W4jgZ7Ow4kNfzizSs1TMydUAD5GHsS2sTe9F2g
yNUIL7y19fdY5v/4e0wi8atDxIAIdLXpDWvkSigdsMGgiaA1S431FHKyb6A9qpQFjTALFIttnCo9
vpy/qW5mvzKIbKsveM1d7xfYAfsc52IDtAknh9gdLShGjcMk5pUq5TfW26DkC1utUD3cWjNmGxGn
Yz1lRP2sp9+4S6rnzHLjlzeATPrYfuQeuiachzL9nEAavti7ar0tqaf2qz6vPCxm2CHtD849wzOl
d69v72X8Q4iixwGIyXp7vzoI2WWtMHBDPrGbCfDFknLV1mmcsvRhIxvxQnlVFMfW2B2sTkgxCVx1
Z7Hon5D9hYYGUoI87cdvnDfdEc4CsYpX0Rs8oCr0bdwClCvy5HZpYjRe7Z7wrjoxhhPzBriGm04P
ovHuBXtZGrS61uAL7wEcazz42057YuieHwc8n7NxtjXMr5tQrrP9XS80LMRR2uSJDi3PZ/AlR2fF
T5yQhRpDqXhWvoTWDHWFFrhiIH4chT0N/grPALhFsr9GWmZ4PxMM0pRjzddMduWjix3hgnCDVjjR
21o5kdP3PzhLcBcFoSNvzcQRnAXNUwiBHipU+7/4pcAt+j8QhOLu5R4y8lpym1xsKetgijl2ccuW
JZrO3x+TKutuG9ABpbetVWb0B39oLlpREMFLXQVxuKQxkZ75+KXpffIJ0jQv/djJSGTlshkxE/Y2
c0xtYGpyO0GMzwc5Jl4CCSf/T7lzwJsHAU1tcT8D1eA3JoeudU/Ou4IAppWxkJd4uTkAaVUbR7ul
xz2TwAjtO1IRePvWjNLToHhMtkA7QUe9ovOah+Ha1OgD4rj5oRo39/UZQ7+1xdDWXwyRbzfZLJyv
RHmgwdBJ8USEsVBaazyyLLI6xBehOc7xr5vKwJdn1+QfOq8HYCoeweeCq2gmFhPLwRShsSY17slv
vo78dd+Llxlr8mTmMhNsWS5UnoqKbQufk2zHkAjZchnsO1bkXOo1DFC06KnC9uriNey2bEdLnpMe
rjFOglZWdA/j1dHvl9LXyjSPR0QQq+wxy3o5QJgeLVL9X1MOR/HoJfqxsXdzHVTfjvILML9gkKhe
xPjNEkcL7Bt6rCHnvOh2ie9/5duWON2wrdtkUsBBcAZ5QIFTO7LhdTYbg65S44Q4cy0cEI7/mip3
rlLcXDE0Cyx9GTVr8EfDVB+jqjVnsV5j/geew0ZQxFFg2syjNLKW7n/eT7Hdly91UV5OpzFlsO7E
d1lM0DRdApQTLRsD59WKs6+2WG9Hnrjs8O+69PwrypAaVlPYPu3XBXZ45OkgeTSzhdzR73E/tdD4
qAk70oHZNdpjWcv2qJKd4ITz1ERu7cs8KyuLpbsZeCxD7edJhv9iSMzS0k8nMDm1XGv7ILQ8aWJE
rengoUUP5hwdfN2a6QzwehpTMP/0LWOqVJyh0n3I1LVRUUntMTs4j84ce8KLBlJc3svK32jArQsH
CjrwPYCGTnWtsfstm4wHnaZumxPgFXWc+THQYV0a7Q5tfOLwiJ6dV2kxbY/qnVY5ZyqP5j7FyuKP
ysAfuztpAdrusRaIbX3rVzugXYG1IULzP/QiklcGoVnwAh5/nos9P2RYmHUM5zXPeX5nHfD6rgEF
oN7qYv5o2XSFfuSKIexKxddlbyRc0OlhGIIPxq93/+A0oBpddKrt8vQEZ6fh0WPpGp8vxROZtS6k
xsIjSnJKCrhh+Gx+nutYGB2H3gvHg22ebpwWzdYI5GbRKuOoPVJ+/dpxrfrb6qn2utGRp6KqE8Ut
OlNYYNFQNVjeaYQxmMtUwQx/Np2s7v3a49K5QZatf6IpLAODYgfmLaCSBQxGcAHXiFKvS9f+0/PL
YvZLg3NmdMXg1bpsnz0NjMcuxOJBqYmWT+q/S103vUFwTtXVrJevkcUo83jBM43kpcFul7km/aS7
EM1qKKF2uyC9xsKPj5ud6h+kK6QjuefRJ44lv18cTGxYjwVFuHG1WxnDUSaSzUVOHroZrR5z0j+Z
Qmaxar3BqjHyIsoJXfwQbWJdpnDfY88/w8FfKRpUUoYkIMm70DV75y6HBUutmhoay4DMZeP11Ja5
Rlo5InUnqFEt7O1djGbrbFYrZUAms6Aq9CI+UF48J1ORLFfSZUIWL7dcOAjlSYz4LWBG6rWUrXeH
mfxZ/BIRaFMKFcu6aeBFDPoP/PpuD0QhBjndM5NXKI8XlfJT+IJG4CgiQVJe6fMaZW0KU2+dlzDn
YS0jL3uEsQGuTnoB4a6FwCXTrzKyO0Na/2A2MAkdDcNe3ILRMmFFJn6hm52sJUUtaXf/9MbOCR0N
uceh82BfNlpy2SPDbRL0ejWI4j5zNHqymxkXafn+PIlN+jTB7/0chrULtOElC4Gv7E9kvDyXJBN4
sARdZyI0diFi7Kp7Sn1AX+zAk4dx2y4zrxdkNNlNXK5MA5q1jr4uUOyEsuoTVvD9JlxWD1yya1tc
4o24ULiN9GfUFdvQhIwtr5ELmxL4WSMOK1yjMP4kTrH9TJfcKwruZSM8jAq/Iahy8JeFER5x5I2m
+zQxOlaCCzoNe/E9hNF3jz7TNHPMB8FBiAWD6Li7CrI9/kOs6DMpvcz7qLDwEuUp/SJqrIhSgCqY
dHyZCQGxykNlbfU9bSgMr3zNQnjC3fM=
`protect end_protected
