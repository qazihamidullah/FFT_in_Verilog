-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vcm2zBhnxJhFQ6U5r72Bi/lday9q4kbjXX3TnclSxJBHmdSVko+eyCbDdsEFDWQ0lnuK3+/9n0O5
D9jKW8ltAgcqldJhgpgS9SFaCyT/PpaIF0yCxSGOCKLTLHZpfCKt0EoSZQFXCy27XDunqgRpyWOX
vB9vN5auCaubkUMuWO933WjK/7d9STOYk2g/CBarDovFFG7KFKdU10CwP9J1BSLrE2b5kNjIW04z
pcaMpmBUAwJkAp+CLUGNizemoI2FwNIsGqqs7J9JciX2LBNEkpMGhsLUgGfSHdmLQ4dsqEMmM/bq
r15e0PtAxqPH6LIROlg5pQK/aozacw9gU6eikA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
OMWwhbVvfhXoxxhyiY5qAGI8N9T1O47lCsLjHFya6ocSuASOaChfHy0sFo8S1p/kklFSRKd+LCoy
0RQuut1dztJOmaDhSb2PoMA2m6Q7rjqdvbRNrHhYGJbe+1F/zUzSKcpQOBqWRjLd2ol4O36dBguQ
BcE46Cwy3pvycnSDpQoh2Js6Qp+botINuQnyrngrFx0vwHkuK9IRYrJ4YvVRlvgvntnhdrSHPr/r
sTbAi/0iRzYxUGja4xQSdMY1eiE6mPnFBEZt6Okr8DXcd72k9iZNCkcmOIB1Pmj/79d0vaz2s6aC
PfzdoTqkiD9xKRgoSuhZQyuigTmtgp3pS+8jYPcr5STRvlxldnSHyr2YQEjhUK2jZbkYdc5EzKno
BuqiIk6lXuR9zEXcLajEb2xzYFBFtB2i1W7s/LCyeHXo6qRFd+wfBkf4NYninEm8Az4KTpjlOfQi
DjP2AQMrxe92P/VeG7Xst1mmLUuvCCT67pzNKXvIEkAQ9sQIIyn6OMLn+D73atv/l1NOXNROaN4w
RFdvKWot8qVia85xMyX4eRGIVlV/81fohdP3UqX9MIBGpYk45gj14RFo4/4JNdM6UWdKJaSQGjoR
W19pZWLtfnabOolD/otnu2A/WgeUoXks6v8bW5nXo9HUKvBU25XxhzJBblFGnI8EyWCXBVw0MYe9
+McjSGLJMG+NZZvRut8L/BqP7OSUvix1GYAwfY5honshhbqnBJjehVYXDKzTirjpy+TY92appROC
FUbFjJMqVSZSfnhMMxFxw5N7pUdkIQIIRYvWgAZafJlbmXCMbQBEC45HnTMySO4pMFMTB5lAqY+M
zCZcl4+sn1zv2QV/fL5U77hnJ/sLL6xMlWKYsaPndjM+idwlWR/QRCykujl0Q+Sj55e9XZCYJRXR
1ey2oOM2DIWF3Et3GDzlBeNvF2PX2D8DZUBYQwGecalCxShpdodEqttv/Dp5hoTVCllpI9vHzHBP
MfWV868Kcr0YyeSMbbzfgkOLHtbCTMHmM265dv0XHBllOrlO0PwhymiuuoiSUVH4OuOQm8ZQQRqy
o1xY8ugudqz0i3SdpmyGCzkaO62alYBhGrWq5iGK0kEpRuxlMQkRn4RqZUXOwW/H6KbN0SpFqeMS
itSafiGDioF8RFh9g4ndPxOUj3hIfRNYP7ZPIHICVOG+joQOmBw9y3F7l3/8l4lGzucxdW96dpX0
n5WTxSj94RHyfGzzrgVwpLC8OOfuDb8BJLopamVnQWwsK4W0RczfTpy3TWzZNFBQoulKEsQJdunM
6SvNBgLWxDzpwMxzU6/OCbw7og4dD8H2yNapfrJxdUEbZYywdkAV2v0rPYC5dOGFFn3F45lcBicb
sCwUw2BJbqZz4EVToYB/TJ1YwCdMyYlN9OQlRXrPG58VjcBE/8CcUSihpGXIIOl8+eEYGGdkqQCf
INXcNGJ5poCDUygDYZSuV7/Qw3rknWhv1sXrmpqo3sdQmKylihAue4TCIzuVOZrs9D5Asv8CZRqI
LLWNCvG8e+AKWKO5Xl7w+4d0XcD/ZS9h1wNi/5fUwGMmP4sYkGxsE7QRo/59HL0lDTrqy746M584
PEc+YLT/xvSw7SC33DS4WiUZpHbrfzIKquyOCYn+gPYsuTiYCmioVKfoIy5DOPLmVW240e8f+ZxK
Z0GugXvrCCvQhWCaDJHbbnsSJAYTOu6RmENJFu57rmZZsOKP7iBksR5s+zjFEz7STh8asT7fmI7C
Rg4k55oned4GFleaBFIHMLzNPCWS4BWleUIhUzgbZcNC+l6/cQ575dHYFe1MrbsQfE9IN2ODqAAZ
qO3K5j7lERvXUOpAbrRLmQpkg5URaDja417j/wdJ+kPCgBzcY/lizDwFXd4GABvLrLPFPHIKT6aG
sX2LadZ+9skeu+SoKSpss6BSYy02FaEIrdNcbCSuayU1hDuVPqRB2LEV7ZPUPuNdISx+/5OumfWQ
YTT/rnJoszjsYWKHESeBZG7aCGiw4jfvaMCLccgCj/vWiC2eYcrkrlZNc2MM47Xmcq6X5uwnU17f
IdlttrucSEbHo+qjdeoQHBjindVRFZEtceND+fSSvX0ImAdOuRey4ME4Ft4S74Da22tqLewL0A+R
69kIaYpeDVPuapkBNYbDeW5DzHQACfoB0doSTW+guqFPDcn5UU6S5Q08kY9ERCFdpYiPsljOvjwj
2JeJ5fYiGCfzJH17nFI/rw06t7FqHZ6tY6vGo6iykE4Wt9OhpkE7igpecG8+6sLOJYOoNMgOwA+f
M/oWRMnJEpC5Xg+s8QWwkgVPdkh2/xBcMrwiFOjUA3oryVBJCDybVRWg4kkthmmnfFpHENpoazPR
Cp45W6AKsgdgtUF+PBZmwzuUHbrb+BQb6FMW9rtwPdCtX/KlJyQE9yuVWdIDPDoUSxuqWNYWHG2c
eN8u8I79i+dEB/ls9Sx5nGHEarTCRxXkN279jNgOtXBMTRTy3jqoQnxkv7DJ9w9VxuInPhhtv1Jh
CAR1U5bShjIDOhI/CghBqRHWR8T4+8Vf0lV7ovbpd9wQJCLtfZsdJkSbqBx7rteeMTzqO4FzIb5C
AywU/gBaFzZcq1oy/8u5sIjjzI6bZ9j0v7H6r0/oQ6IBX6LhiJmvbYF4TJngD8xHNV6ibH2gNWSI
+qmH7nSeHDEWkO/0n+WGXQCGN7H7mJabQnnIiV70yPoRTCIu1rESoDUl6wXZqzvqt+/Ajk2pW+LY
S/Privo/agJOxCet4uDPW1BRhYIyVJXApYZEnO0RYatpxOj0ZMZ0P6a3RCvfQwkMID564eqXZcDI
2Hsy0cUwjg8JvI8F68Z5ERQvwdlTha18GAzqwvIhbYDs5hA41X0fFn4auMT1Lrw1o4QViFeHHQ7Q
vrIX5mxtx+cUZYwAScnPIe+nWNY2bIbaVLsYptXq3SCulOmp1cHhumlaP4DNIDosifOOBAWJQVoq
xO6952pRBWaD3GoFyf7obYib/E4EjtuMuDHnPvoNgIzU6rI2rJPoAz1ULczIJ3y3iDnXLRaiwAxM
+20dHJf41lvDbJjISxRM06EQ/dyOg5L5VsM8d42OZoaE4UFI6BZRvsmk8KPmySWXED1Z0xGo54Yt
Jbe509lkom/rMDH5DrqG1FjC7R5YiskWAzdQvleohgksjcT8Wv7kNzTcsUIgMYYfXNTkOMEo3rmQ
SP3RAvltiXky4DcDt1AeOV8I3T+XWCi0sLFPmaOvnafp6PR8Feayzv9VwJEkXjNpPqTmnqTD84+r
Q54AzkKSBjBsKnH1NcldIlkY47LarGuHb3Agr20PE7FEgL/p2aQ4ndT7bPm68siw8ow/EbdfRVVX
Q5NtWZVqYUNpVET6uT/r+bBix4oxlFndTb/TZfY6mdgYFBNycsEfsWHBLclj3qXbsq6mmdYlGhVu
R2XyJmMrF5oKDQTL0jkd34UpOzEacV5Xg/sVOI4GQAgRMSuCZ/0Ntfi5PFDpy9o+tOPJOY7Ye1aw
5wm+u97BDi692Qv0Q510rN84OGll3POD2UPmrHvxJReYHYXRNBwDFzRh6VCUz5cM7sY69J2T38xp
G/jAD4DKGR3yEekmUekrhmjP9lrCY7mW1OxafnUE+jTwprpP4nd0urtFtEDMVuwPxDjMoc4pVnQh
spKU7wY2YzkkQCFq9s9GhR9cEpSy5GBrb7HoZAPKEKmcmgbL6BTStZq363C65oPAM6vAT2STu3wP
4MUbVKiT6yUYA8A5lGC7x79PabaCoajLrK3A/yRPzPW3ls88GfYGIqeiz9IcHnDtGY1MSYDC38ll
Ml/Zd1LH+dMuvBkUC/LhXHrSkdPN6/+DX8z0ZjtxNYFFMY/N3RzuuonN48xWHv6CyGAjdIYRvOeP
bVEcRkiWdSt+tuoQUE0Ep0PxpsWXkxL58AzwPRzvrpy9oZO8ANmB9p7oBnVahqusXwdYLqCf4e0b
IhcV+OYmN+H3ISA53ssJjVZ6Zc3tYPmn/PdVphGAHYR9QZ7i6clZYtqT0L6+YcHTKyrFWxfgmtMt
k1nFsqXv/rymkr3mvZVpy3klWBq/XjWTZFUVXzDv2LZ+cZZ/Cg7uasXtwgIu/oKR9WbkMxv/88fH
KrBRLU0Q8dzHLMSrEJ2KgFUAGDvR+0/NNg3k8tjWtryr64qyKHs2PTfdzP7eJl1pPlxr4FxMO4bW
bpL4PfskytLaopBq/hs0IAxmd2fAsRV9OHZ64WTwD1dDE0kWuf+5nZPKfI8cnTZm7XCExs7kQ8F+
4HZLXT35eS7b2QpgNM8yuK6lIks973H7owIHA9PtIXfElkT8PQ1hztHNWPCF2qwxW80iqVPq/aZB
V5hMU/zHikp8oRutXZhb1YQW6CuRiDXm1ow2ouBB4sxXewIP08x5masrZ22gUbk5u4sf2Mv7tE4A
Z+tE1suARpZn3Q0ymWtWcYEqngG5dk0kA8jcHLiV3ZJqtIhXjBTj1c7e1QnOqpL1EVEvmyA6UYCo
fri2RElJxWEb34i6Q/xJb+YMXdM8j3WT3rtWS4SS3vHdtI6g5GVrbYyaGziWl6tJ2R0QOUTF1Dqx
bpwprdEoNSVq5cjGR2IwgTH5BAVAuSQ2MVWbvKvsnbI9yFBVowWnoUl9QCS5LwgBZDmH0xEYnH+0
RuJSYLRsmCMDyScRdXPgeCbuDuGLtUnnqoebCXBFo6jLcJ4tF+6JAn4IWq0R1UbDRRpDBFLL2XbL
7sTtp49L6tFd6D0VETxqfYM2TBEjlau1bpaE+tBI5l1WT3A/l0+X/6OgGNiBwycbQairk2Wk4as4
W/yRm0Fh2SxvDnnXxJ5qD0HmZWJ8ifmRTmojB7nS/XR0I7ly0GB7gNOfTm9KD2UG4EW8ZiieeXwV
pukL4WGN025ha797el83+Gnmv8DWNgNO0WQPGIh8tjfEJiTSj0ifL+83IBX4x3xin1dt2G2EWonn
X00BbfdVPuTAfsoyT3ZWvnynUO1lyb/Ywf23sF2mXjXoXhIu8fmF/bhMM7F0IRY9J8t/8FH/OTbQ
hxqAxQxpWOe9pEKffFaXotGVeXK4+HRAb8QGXmbrnr50elGtz/51ZRP1pc1TMtY1tI55yCbnu06q
EiNE9yGj7QmXeRRUiaHJHg9TGJlS81xCpdLLTKuhT+wem2QBgJZvdrYkZ09tmo/20LDMBBVRQQOk
hcixR22R1LNzwVe/BddK2nJ1FnEpURZQNyxexDVa3ksQUnrrgb6/WQzac2etpST3gNdUzruo9ptY
kyT1J4HTEM/Aj6gJ9tc9jIarf15TkHAyj/sJxK41SXmsPCzoM7bjHODYN4X4ljcx5JCZK/a/HIEw
BqKNFGP/dGCnVbBbEDcP4uzpItlRufgEewPmi4a7lgjVuU6esfEyDY6p4gTPFVF0P+THFQhS8GFG
y/w8th1tiiXQGkPrtWExWXhH9FPrNvrS9i6ct+dVKOr7JtBxEGMp46Qil3BwR8WA5hBseEiLrzis
M2F+bj0rMT+ZE8XI8VKVeT9n38Kdd3/fW5942Yuoi+Onrp755W4CxYZVJUbNrT8y/BkUD/mGBrE2
GUf7fyHzW59mwasKx5XLwFmQF9lSbEEoTmmq5iEHAq4SP2/LltKwgc7Qn6Xi60YxNdg1GtPJKkwQ
I4N9gFlEfD0jSyGiW8mYJS+UJmy8SM1CzSwbelkRHqhLTLE3nB2dwz76xhAPvvBthEsOrFEJ7tpm
RRWsZIdj/n/kP6hfHw==
`protect end_protected
