-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
yJJTrc51U5Z3EVxXo3+NIzL3JZv3EK2SLQMqm2aXGd5B2tcT4sROgKYLH+uk+jlerlZTLtOD3HLv
U4nTgpub6tw9NaqKDbRUSz013Yz8F7EmlV3FS1GdpqLgDpRtX1Xszfn2Cq/PzTGdJNSFOTYSC3Lj
G0HbY9hmp9EI0S/ENtiPsNvO02hLdVji9layagieIwExQ1uw9Pv/okaj9hdDCzflMMj6pBYrOI2/
6tvC7zN7/yR9kASfPFgYa6WwVIx+onLDpAMSVkKvCjQ6Knu6nJYdh3tee8D6QtElv32iDGJFHzBT
AngT1aaGLpAsviIR2yoNpy4H2/TyfLdTjfQp3w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1728)
`protect data_block
OwSzUzUKCtqN5nY4oxBh5kkFFuAK+H5vwIXlYOZWXMtBcYE5fTKfoslcg0ttcLlQNDHTbKRhSAEy
WWPMJvRVB1wWc6R23oIogh/iRjywxAH4Ne1C3pXlGyPeJzujcmcv2RBQVhN6n1tDqWC4iYkI7p8m
P34MNSggFiH5gR9g969zSbeYqqVxgNjG4udhTYyuSIxw5sI6LaFFjTQHh4tWuwjQfnwZYPvpn0cT
iSwy+cOr8Bq7li14GmgE/i8XntZwRs+8xpUDb7kYOPLBy1oxzsoGRKcsBEtMP4YVBAFipu9jutYY
hry1HL5yWUreenJcQ9I1EfzzHJSdhy6e6zXW9mnAdsGaPuFlgNsU9hVENgwkNG7e8Q40qg011QqF
y+PCCxa8JBy9mIONKRY8zEsuUV8fFgCDwc1hPUWYUURYVIhNkDsI4582Qbzpd+/D73n4pE9aED/G
uuiwKyeG1+/506nfWv7K7xhMepoqGH3KCHevOQBp5KvfNmBjlNdycTqWJsBJUR63Q18zXDnlaPoJ
d3wxwrGoYGMS+bhmeCzZYlJDSq1AWZ2oC0+kjr8bBeWaIw3eZwXwHiJRCwOth/WkTVKDqoLpIuyu
W6AK5AwnvDSsM4WZhS85PwqTfWC9QByCqYzvRgnF+o1OO3OX9brKgM4BpaN0ulx3u1XLT1OkSRlt
8AIW13fFPYl6uP4rGLzooUFYtYOdRUbZi/7ambuvUHDsoX4klMQjxkIcIhX7m3UmpnfP4lj+/S0h
KI+LNbQ88xiZHfzsD+E7RHmnUFHv1RuixJxNNIjcjd6nVc2qqY468g/aG/z1z71cuOAxOXULcH8S
xhM9GqUZGSR9BxPE5mnU/TlCt/p19+qjIP3v7eQsvG5hYYl/+2xKUqAbQsi8PGnUDZQPYsea3hvQ
exu8xFXgJ4h3lJ6Hs5BEb8IArpMK7K5WOJ9wrmUyAKd+V3lBkwM6Wd8xsVtvIZqkBT45on4uwmH5
K61q3if2Jjo61puehM+lYOwZ/g/lhBSlHjnRPihYROKu3m/Ndet1jTHjbqlHKecYvhrQXPtx0Inm
HyqEm8KvN9WEaZIBMk8OlEF72LL1rmQc5ZTLSYdwJ70Ensw8gv1mxbvmKcJNuaBndyOVE3l8ol5k
q/GUZcgT+3k3yxPihCaM+PZ9dWEeCtOAoM3WJr2eel7bxuAbMX65xS+uIIZ7zdB5olgRjxZMTkm8
ZSGxs2sl7MOZvEsflPNdlQJk1DBs9aCyQ2R9QU6SPT1J5tY7PuCTumljW/5EWX8dSjng/5mGQPUg
RrX1t8bzTS/gEMxz5nsqnF8CRtwjebRYESwlXnsfCrji45gjCCZBHHZDKeU/PZGuvC7nR5yvnlAG
NtdHJ4LU/3KvfY6/5EkZUitiOJlMbdZnkLZsRwsA9ETHqyrLo62mWDXN+eK1jw0LCWwZvU072Ae7
h2XOZEshBvi2X7SJ6D+he6NYCjxa64B7gMHycslb7OURyAKfetdpRjQGOb9t2giVkr9NgaHiKVCW
8MG+zftYJDi17JvTebzEvoq/CiIJs0SJiEAeP+AcDem0Rpn5CqwJWA8zDrXGLm0zwKnt8tTpSvgM
tRCXOu03v9RLOq3h420j/xG1BevDs66JTzaPIhKXyrBhXP/s71eWf8xyK4HOWLxnhYghs5+V8o5x
OvZhIijs0nUEZrMK0aJNSm9W2n3Gh6N35H39UGPo+/B4QWzhAAecdgGjNe/kjV8b5jDN/ReW3TU9
FLjSBdvCMr3hpFFWdpLqA7fXpV+sBln9j9m4dy7thQrmg1UbNzjeu4BhUz4B0S9V02bo8aqKSskW
O8GQGBu94DNwYs8jsxfBoTRKFgqnI0OdyhmhR1QRZSPfB0zUKq2l25O19VgHhjeSgjsQrUKlCVWF
etS/wsjir7GRurCHUd3hsQ/46jjLHjddetnY6TMU/6aeUJ8eRid9dVvJLu1FuYqAk2/lcdj38ZPY
BDq53HVXtcL8l2+JN77esTzmTcjCTaJeNVQ/JcGusQAWATYQ7/G1KXxUzj8EBWfwIXB0j5ASzDCz
qgPZGLxpXPFpeK1r36SPYD6IXYAiVEi7v7O2+LquGXq1eYgXwPVykns+lFmhSqrsB/QEUvYbRxpI
3y/yhHuXFE8eyndvy2ywN+vEnyx7OXIWemLcIGZ+Ui4+7+EYCTaWxCVQSfC2OCI2MDEaeitmFj2F
A6GtiPJHHX1/F9gVdFYvqXrEDEcDYgPvoy8g+lAtk+izaEcqEZAITcEJHV7QZkGC0ZaiIOeAlLMB
NPUxEkpGCpWbjymnpMrY+jkN
`protect end_protected
