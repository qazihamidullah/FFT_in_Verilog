-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bINlcho4dX7FRnfAsBMdv0wARsdOYZQ0PYMNXyQquMagmtkUyitzFCy7HiTIg4wX+wGQo51XC/Ge
omwK+1ug0fze0mzsNwn3ljikc2GLnaTeqdPTKzsOZ4MCPZ38rcUJzqecRPlFFRsHgZLclLqXp/Rx
3bQ4cNlum2Wx8B+ceqADvXfpl996ZZyT489lBIIjvHwVlLMxz4YmdT0a9E6enNQuDVUpIpsvznCj
W8y6UpTFCKhwT6ZKnp/h6iw2yE8MB7ID6E/sFRdgVu/13+4tpsv+AZFLcpMglrjkUE1axR9rt2Hc
aqiAZzGWDztT5BnohYyPWviu6Hy0ziAP2JtM/A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4528)
`protect data_block
59AWtCkyRg2lT+1e+0Tq7eEuhu5E6qV4kLetCXOZBdOUXRdZTuvLoZGFl+AxDZwA85l5dpEcEyI1
Eevk18BdaECjJzpH7cW8/b3WlUQ4SN95WleodX61rZcijiwQ/lTnHHEsR9owx1eJwjj66ZC4MZ3w
gIvbQRAmqOB50txeoNRcY9IDNzFCz2pfzJElpkzQ8oVmKLA51Py6Qyt+WF/aSa27kRQ1sfQL3KRl
++E0SjduQX9iWtx5nkruHcjWI709IcrAGuUfwEe7Cu/+441hA0JBKaMd7NZMzcdXLN9bGqSr4GQ+
Ygh1yOPqFdQHvVx+12muKG1WYgzWUctlt3p5Qnkt8YBjTFuDTLmciNmzyC+lskUU/gCs1GG41Q9l
8zBwwUNhjeykJnsQnUv+NzhO5Nvz2sP7gmogoOAV57MS1ZfC2Fleegvzb9MjoTAiPQjLDmsmZMZU
YcIlcWP56gQ4gOk2AP54AOgs0zKHS8g0/d/6Z5CJoKVr7qAXQiphs4YmeJREnGRnpcBs4NsXU2kR
TlLrox392uKmv3qDlI40T8l559LFj4X0U0xf4yQHHQFOGinFL960vSUyqzPmB02X1bIPDMbOMI2z
OmCyyfUsRTsIOyn5D3sL9q4X55GD8JihVlYwnsGCUQzuVALzjWQoxrCGdSGtNKgv9AxSZKn/FQ7Y
X9P+KFQkUOCxTm1D93EmmobsyyL+kfYtnDnVvaAOQaFGHSOvlp6NmLQvhmHp6PcdIqcnQEqhz9wn
LGH6cGnKbSUNaT0odS3BUnucKxH8YLPxH+PY4qYG1d/cYf7pR6Ou1W+hF+euDUfeGQU9BhZYr6M7
M09qRfo1RqfMIOQRRqEU/qN0pYrKzUEUr2zcoGFH8Y1BRNR1BcP/19zTgYYEO9qkXJQVbVXkfh/o
czmLbra+je/tKweebnZGmGK6qhKps1ocbs8wzWZLaRunJnShqjaxonFvHPYdADkMM64Je79Xh4Tk
vSseFH0YswAVR1BemQdcdm3DgV+7p6FxSgqGBjm588pn/B5w0KIbfFQzA2dodtiwMUpmMpoLxqw3
aiV46k1Y/icObg5C/lzdJVm9aMesiIzHCuJq2FMRvY16XmY//Xh7kgwhjYatCkQs5K7VgkjNRcj1
hMKoQX7UurFgBy7RSrvrDUdagDS8O4uCREGoIfgyr9rX1iMjLDfwQUagd7wTVzILvZhRMnlMmZcP
pcbAKk7uXH2iVX63LY3ujxQqOC33BdfzsI7rwmIX/XPT2tgghxTtD4v4ZXgpbPiZ2FzpLTJdhEwI
Zsy8/4d1fi5ozgtbrYe0u12QuWNPe6I7SmwgzrJjmXMFWg2r+5tjFu7EuhFlQHZBDtettbehnH75
DAEjUEXzuAQVXj8Ksx8aBhiyIiiayw1K7VuCkqBJhYkN1Y5UIN3akxNShHXRDNNAM/X+rv/2jt1r
3wYaNHjPfB0oZmUWuEXZyIknS85G6qEIHuiRnC/VdzxPbc5jW/0GuGL+9L8sMx6CrdT076baORQ8
2FZ5+VI/8bRMfLkTFT1m+8t0yiP1Ji56D6zC3yG9TpeIznZQdx6aPgO25jF0uxxVpLT/AQ6dEMXo
vUtCKZeruPNPD6P4SGcVL2EOgHPas+SJEtWgVvl3a2EWqXTzPY70EJFyJdy7JkgiTNVzbVTPoDtd
OELh/Kws8Oi7ju8kSsi6uiNHyr5zh6JwmP23LKI03D0p3kC8pFGaj8CACQkfW6E+1uegL8PFlrpI
qjdDfX0aEUvlfXvSdlOrpFxK7WOxX+5Iut/8UbofCwJ4hf5EHdFnkR0ZSgNyoKooXjTuv8SzB5ov
q48y07EFy8PG0+Q/oiGYld2+kzJ6LRueESRrLVMJXOWN5reFmzeaIOKTBMy2MWExZHlWeLn+IYyz
OT00AnA7EnRBg6nJr1gBPCjQf6PlsoGBmzfqe8PPOJjO2osA5V7ywbWO2YLPB2D65O7TNOmMkJkp
cZsT+pS0Y3SavQS5KbG7D83m9Q/B/TjYfFL21GmHU/uLiIkGp7splpX3muiVt5EquaNg23JzRyZ4
HdPZ2AVgBD6BX2UyZpb0MN72iBOr6WYPhW8ngsb+04IA/5og3um+XrcUYd/TGsDMDUFccsmtgyFQ
piMF4u/yVrwEYCOFKprqhqStc2bG4k9cK5WMvHCtIS3eo44nrKMuX3NY3mc1rEsKb0+mzjtgqTVs
WiBVdKxMgj2Gemf0FfFURE/eIT4VbVqwrBEX4pz3Scr8Ig8jYLZ/oOXjW9hHawl0moaPtiM8Hd3R
xnZiivkimmJ3vc6KCW6cA0OHKxhZGbXZ7RxSGVliDp/9fJ+pUDe8XTdDp/a/s4G0iPMh0h+5Z06W
rWSJWrvPNO/iGyIFwhRPvP7ETt2kJvfUAob8W0dYI7t3lWxPrBhO4Lp+HtSy+U16DU1aShpYqBha
kiE6F1YtuQ3xn9sypy3KJRQIlUKGJEcJmX8vANavnVoucD6/X0Tp+Cc8Dp+4Matq0et/cJVHQmbo
Um3SqqrCSgtIu6hBj79+7thmvPuukxXI0X8LD3FJTJTMwD475ZcTB5plj8JzjQ6GPoVqYdmbv31G
kG+HtgOXVOg35keCgs9vxTHzwDZmUcD+p6fq/o/9jP97zHVqQuIBzA0uxVhMlYaOA0Z1ZpWd5rcG
10x7S9/6UMnUrDXt0+jvZ46PIqIjotqZqI3k7b4dgzEXiGy2K8s7OUCuWLEAtxrTVtjh9XSXKM/N
5pGHuJjOExNSAsfvT74cr6LICG/RxgMNp7Y1F5LVmZxiqU0ki8AnXRu4wjl1N//rMBSopnKYi7Sf
M6YK7qUB847/b8O0nrhQ96iS7JF72+dlB0aISNZyWsRaoZZqC2IGa38SPh4Vm4xvpXFtfWDiJJ99
oY5oslprVWy8wn8fc5UF8T9Mclyw8kWm56IJc270Qj4g3ZoXaxemsI6CDgnS0uIDwIRdPL6jmWak
rwA6fXAJ4wj9Ejzv2iGqJRxne1n2/BvomjLpSIjYQR6osXJXYW90dTQuajoq5C8b9xOAuDsWfTBq
GY0CdGZEGXerBkNuPS2xjS6br/Nz7dlSSWVAmraP96+MCHrc2UmJkzqfzgXCOcu+8yJOvF87aCLD
oRSD4V1CokCb9iy2rUyUG//cRgCTZUANLdL27Katy3hq68iHE2IKRzJfl+0HTUH0mKxCqUiGUrlh
Nr7dBK3Z8zQkbD0EGQC7CeYpfCW6xsoGNlGFr3acmIXMev7ORwaOnDBUMA8NMtXnxKhmWDHYCWS6
vZ1jt6HxSLJYKnl4xJAcBXCC6jv/TFGHJhA+XAB7c5ZzAmsYA9u+51X7F1oaOIWgX+cqXOy0RObO
YIC6aUSwBIQ4OVRxBJh+zHKqPkodOFn7nsC5xC2+zTfpRnNreHRZ2GyopxfqT062jJSLwwfwaEDs
abtRGNrmKrZsnms4I4IiDz/r03CaYDw5MwUW7/JiykYzEp9zpRCkjyr5HKKrdnThW880TgBMiBYp
UE68fe97WUf4GeXN6X1MXDwB8W9fcXUsCDZo7xYSppmcqfCwvc/CP+/g5GekujBo5fEVgdkdv5Tn
vxFIYC6c3YB8m991zPv6juKUEBMKGfTFzDSO1oevBEg8XFGGWg2fj6i1in+XgdACAPk2p7C5Ue49
tSi2np4DRW1hCbAwdqGXPkRgizAOo3GEG8EDm++CDzgwlshpPVYtMremKXDFIHeB0vqG6NClEn68
l6lbrkgctKTKuxjRZFqBCDQb1gpMOXOd6ZBEeNfXC1eqsczjVgNANw8GMsro5BIAGwOR0sB7sYyl
bVDfWZm0G3AmcXHxfdIaNumlpLpnqS2P6XKEJ3XKB1+Axs5zLIJvnLx9UBukTJwXdDsXcFdtLvxu
2VigCl3MLuvxja9Ns0PViNlLYLDRntUNXBmP6WtX72wPSy5dE61hgd4pWT9ncxw59y/gXF448+01
6mUFNcbWbAUIk2lsm23YmVXMB5CfFV/1aTu0aDWGFhmgADBh/WiN6sl1ZAkn1oQ6gemp94ALBseh
hCRxIVSZhTCATKwj+aNL7B2+vLUUQtLe93cIxfPjhm+ZhGooNWBLQfU4eAyXqcgO9ZGMg1loz9t0
FhbKkZ5xVSx857FL0L9d/LjtjwqMbVzn8NlMHk3vly8AMZUFIv5kPd3W5VyFhsgTJ7FQn5jmK1Mr
l6pqtjoLjlK7VBOQdSajqLGr8J3cxxs8AQ0zaWN7XjSuxKv+wcplzN1O9XFyEoOx74UTKUREskRi
uav5IfL9+Ri0YToGQKFjaEhS5hKtebeDZYDXEJdUaSfXRKNgUPYjWHDQRKijfEDwY06NUBlbtiRd
Ar5KzyAtBHSbOblmJ3Uae3GOSrelTz8rYYIZ4/Mxz7Lq647sGJc3OnnsHrYz0e/uvM1ZhliuVQUf
bYkwJolXrCgpRcqhCKycQRfgc4LvxbBTiuIuBHnEHPurJONW5YOAfRx1tE2FMbWmznthfnKddRy8
g1Bnwn7hoJYhTKQ45ZnylueKKNukqA19B4k4JCQy57uvFnM4iqS4U2/kee9IInGzkXWiEcA/5A2D
HwnZIe3DVgRihgQWwMEfnImBodlRzePUvZSWqvdb9U4A0xzFaZfgFQGPrI0lr0dN3wbe2ksFik2x
5dnj0fAPb4lHz2AxJyyPDgY6UBoWoSkEA+Pu6iE80EyHTsbpAt4khGQrKT/qJoL1Yp9Bor/J6v7e
zvBCUJcj4QrsKnpAHwgI6FoLPpoy/Kh1Zh48d4ROwjBgYUzLSLQZRp3Q4YdnrcGWae4HD0SJz95g
QUCg5cXfOIbKnUV4oxLx7AlhZ3FbXIkpbDIbQF75pqksdpiUUoa2j2Ge+2+hVAkK7WwLvluvplOK
TgoO2lUouRQZmEjaEwwa11u0n2/iXtIOlp04DOGPTD3X7Os1MRxUWiipFSFUb/+Fs5ekNR+7dK3i
AWka4iKojgHgOmEUKCMHdXErbeEu/gWgCHh7RtU70X9RVMuF3zBYb4EuuNlM5ehdcIyiJfFXB68F
VKjNgc6WH3XA5lkM73PhU/O9WWrRZssXW8giEkX1IlO0g6THiUiM5ROxf12ZZ8P3ZmqmGIvHocaQ
fXSs64P0KOVkyyq2EYsIOqmoq06V3CgYRxfbioTbXFOhwlnhHTjppDX0l4dqFlhQRRulCtbl6L4d
zpsVAr9HWn/cJy2qECHJuA3qrgpI6ahkQIs9+H67Kl2nePrSNnuo7wWetnhr1XEsZBp+YQzEWtSw
oOBUjmvmY7heTfV7wIyKHdZw9vNCyihoquqOON2pXHzrzTSh6ZLsDGZl0krO8RDuz90xQv8Vukzq
Dd5YOmX/e+K3p3AlmNbWeNSuCWo5+nFQmZt/ibDEQ8ftvWRA9Q8FkvucKTIHdzni8fNYTR5Iu/zk
+TwsGowkrYzoRFvz7B2yiuSc9U5L9G2ZYop1cN8u3GARXhsKpp871V0ZSALHH8j9VOi4M/vhufK2
h8EMqKY5/c8Ff6tqPQdOMOiqIl6zyyOehd8/G8RZZjflwup2+it3jH7iD9W7MOyiJrrWW+L7M/h4
xMF/S+icD0jrGcKI2FlRzaL09+6OfKSAdQsyiH/7v28DUqY/EpeACNDQIhmYUTD1Va2WThQxvxKQ
CiKIrBtiTZbRh4+HQXqpgf/PrFVWCfrYQT0u8DQDndpRjz4d4WRFa6PaWgLXg+mSd0os57xFVHOe
g4QyRXFf2Q8QDF0DQA8WiNQxDU7AFWtNVtzp3WfXE+gv4oaHTFr06FeGgrYM/yUGva2l8mL+U3TY
hfUUcPEyKfi7CljUSJp6fonWr94hc3N5c8m7NtktLCV2J4ljnFH/ixzotrnMjdlsT7AxDJjgZj7j
aAcHj+r7LFsFRt8QQmO31s17+MlNEJ7FSwjKoZLN69YYx5Xezw6q1kp5i0kOoNyZD0Vj9MSCksFD
Z2uVicJZAYcTkjDIiI8Ewvb+H1fJ2tSh5uQs5P2cgsR7fy/fxkOc3EJz8UDJW6HfVKWZl/j7SXV1
wo3Y2ccbmbKQjpkXLCeiXOyJlCMuSmwPgg==
`protect end_protected
