-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
X/+B4eQ8AGXvIHtBZH7lwjz7Oi6Ixfhl2XHjerf1J438yujf+wUVDhDJs2Xq49jjiD8W8LgRin9M
w4F7+y1H1xl7BAzRfHkXCwGhwR88UCS7SNCAg+H526wcXfqu0GIyPELUkvyc/BmJX7Isw/6qxvJl
pS6ZuX8X+jzAH+wjf63L5juqVeEs2ba9sI2wo5uyudbRW3yi3yTFs2Z3TcaBZvze/p8WInCQH76u
sPFEG9TKfP+ec0ZEnsZihzhI8/gVHzxYqa8hIDtKOoUZtm1oovPV0N9JXs7+J0v8QpEjXF22f68J
ERSnCUA7ZAuYPba4PprtRdViDd7kL0jRKI42dQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7936)
`protect data_block
AzHQVfpjAyxJstUU7NzprK5oaiDB0KYhsLVVTAcjC4m9WutwX3h0h5Klzcg6J89XlLhuZHiG1zus
4I7RAO+l4SXcmghqoUPJAuQQuVrGC6qr/QlG4pnwnuHgEVACH6iGOSgkgWuyp9514fHEu0PgVMXV
JjNpehmxpwQEYgr/5WTFofPIOKPk9iwPyCVU2PGuGKgBD46jEAoFt3Ygvtr7XktXZAWLCY/v+0Uh
6hzO3Eggu3I4KDq2uH4X77k1eJUY6jOAWY6LG2Yj1dnSJ78/Y7FnWvTsuK2gu7b2XxpPEc02fFwe
wtKindNE3wdJnR5FEX5sQSUkfZcFIi5YJoCtxVBKcCz9szh+/JsU9v6jmlO+T5hIz2QtX2YqrL3h
CXNUpM10VUEgxraFlkLr9YHTEo5Lo9C6UiJBeHrbcsWs9XgqkhqC+opvUB8F1w/JyTRsmxIoWk3Z
ihyy9oQc40dC5f5vFjP94TtmvzQ0MvMpOg2GpR5pBO8LRb+GjaHPhtTLbyjU/qbnOGDUr++gcDkU
psuN1DsFsGsOqOXnAUpqby2zofQI1wD29CJk0cQxO9qp6RIj4JEbA7ijvRF5lnsVODEuqhD7mMyC
UJPz9PWcwAP5jjcmoAN4bdKqJyz+rg2qjuQIGDNY+S4QxFY8/QWluPTXOycaVx6N/n/041P4O72I
eltkS4Hdeza5UrO/9CvL8ePf7QmkHbKzI5QMbJdpw+NBVKn8agfhfk1Y5XThiahre1SOdiUVDHhL
mpNl8HrJ0caRsbpu0U90d+dr6eD4tOpssmDFj5zSarPrmTw+90kAVVeQNlcSrW3oGQZur5mK5smE
aS73ucSAnLnAod4yP2Hw7Yq+BZKSvWqH9cv1lsAyc0WXMztOFHsj1oBNNtqiGmbP/hkPHCF6nVNj
nuOjtOIviB1aqzCryx5opTJJxV/RpPXT6M1OGxKUa3X4O8GVyu7sQylLDpMcVcegq0Ux0jLUN9ek
1H23eBw5nAg5GbYUzrmonFA0bu3jwskebPZfC66oc7jkGCOiOLUUQ8HFb9WxuDa1/TaBR2J/iJQ8
GO5NUDpEFPXqJLSOL+Mp5OhdTA5QIQn5/2yhwJJFhS9X4Yb2a+KOpX4A1ECyH4XYW9hWCuIlxfYX
rLHBA0ye1CjBEez1aku6PlI8RBITu+waaoeNQsS9et7pdOp6mgQixxl7lE0///AiG7/tf+scwhPU
ybpQlSjJmFHZkwpwwvUxIEYvOuODGFVKA9EEtERgLKsy+YwqFrXwQ7bslIg4PUB6Vr9y/9VULGFx
2kOgECSpllge0a6bjp6J7LxpAjczi3T0qcySt8BgtIQf8eDhBR8SSIVlS4CvQXVQjmKGLpAjo1Ry
buCzi/IUg29bipqF7vcsnsevz6TKloz2Z411C5h1kjZY5Cpt8eqhpWwWFlaGQuSyA3FEmdo0T42d
p4/KnuHU50RuTTTgi1S81V8DAdLUNeWgXrSwSvJ0onYZ+80zdw1B8z22/mUVbG7ii6qrz0/otgxW
XO7Pxr4Z2ToAl1nPz4PdPnMnsW7wdcrEARsYaGlnhTag1fsph04hZrTxzTWmd4VS2QUCTyiGcfad
fFy9bvh8uz/B9+s02DKamRKY17LkRMIIvTIQBErOfzO2OtUFSiWhOBqc2izqMndtLxC2kFyfp3wY
wlzKaw/von0R57XA1MYSzuRPsG19ur2ceN+26ceZNi1ih9uKEEsHvj3aRBYSUDj7nZ5P1verkr0S
asPYYkXHIH2FdkuEN0tvVr7N5wbYFysEBSNaDFlVqZ8htqeZXjOF0QjBW4nkAV9N5zH+isARj/Ha
0BXN2obhKOJFJKPKTCoiukYE2+AX00Y5pmoLyKVUPQF8fxqv2kO/7FBFgl9wAhBmEvEjd6/XQ2Vt
k3pKALU0y9tR1RHamX6uVFqEwDMp6AZyBhRXWxga9ggdP5OEL4IQHoEuzPB8fyFi67DCM67aPEgr
gpyrtPgUjhYnnwZx6MIKoZw36UZeUqaelL01MfeZWSXYptemwlcWASsS3r5+APRVhMAMcnweM9JN
Flr3EwH1Ecn7GBxMb1vkk/udLpBaI8asyjW1Gvr0Oh5CaELRKEL8gN83eZWio//xqYdDsgM2De6w
UyJs8UlgjIHksuQQtEi2nB0rl3XVYTNl5Y40VnxFJmPhwz+Yo198v6vhotMlnrvtfpggImacYUzM
hiumuqxNRfjadDCgHft+k4ArRcFjDqqoiZAxFUv4Nrn82uAD3RkzC5LfL3p6MT16qdE2wNSHtp2X
lbQUMPcHfzBSLRCCawtTKddV37qwO637zQNG1+nhjmOef9DDWlzGCCoq1q9xXTwmaJn4VOUXvGZb
C8ALssoNswMr5tvPFmrph9XhOea2Rut9KNCKkystqicx3a9JxCtV0KFO8JNzpVZ6SkSjlI3+IAC5
16pki5XZSq/GJF4FdrshvTwCsHetwpI12zGUAkM3LEkx6+P8Y8idgiCYbZs7jRKZmmqDrEfsDeUN
37pOZ8+viJ7kH0WIx+HkV0OA/GfUw8ooVQbMz6WGVkOlglgLs1DVknYiGR5OKkl/UbRry2GFQ/N2
06KfP+9aiqJyRONAVaqRjf243aSvVUVfaTO0xbQn7iCtzIYoQuWod3tSqJerkIOMnnYMrZuIvfIU
XBCnTrL8oqRclJ45qgo3rfJ+U5P9hOCxE4sNxpGqbZhpX15Wuo5w+g5Cc3heD4OOJ92zqJS/GBhK
vzxiJ9zHkwYa0wQuWLoShL0+e+BVhO2nxrg1mgSCkw831T2+xPF2fmZk98atw1LxL9vUwxb8k7et
K9+i2iJYsCtIo+o0tZacq9xXm+tJ2e0yJNvixZnRel2wev83i74tJNGzx35qaAETUrknTnSgzO8u
qfJUQsZpcfNznpDPE1xv3UTHlmdbSVC46f4bI/fPCcHldOG8f2O7hrBKkRJhQE0tgJpTREBHc8o5
h6rZ4BefEVCgVUTAoSEtY8l002T9zLqLDkraYDtYs9NFULhsKfPvjZLXSthAEI6Ko3GzJ9/iuRX7
VzmKqqLlFmuB7AGE1HIheSziLbkYV7V+k2st/I1qPtbH6NuSQcp/efxGa7Ku9hFU+x8ubWtSETNV
Y2tChx3J37zN8l1Jj+L6ipCOcDOdwskgAbj2I6j08lsgkEj3JemfVWSAqP0wrM/LTRT6IFWAR1AS
bomA5CFxUcoLiQMXqAO+1ayB0EbTAHmaAwq8UmWC4wBxMKdbyJagVA9nER7DnLfsPBypkycNMvUl
SyFDi2eiTjOFCMdSa34CPUoh588sJvFTqlwM/PdYfs/Fkkp5N7IVWsvl+scGktnNraOgZmUMu0F9
XlgAh2JjTwwTiypGVsnGtNoDpeVmhTNdg1vNK/G0ggdH+lRjTa5Wxijq3IWhSo4eJ3iCsZLQEujl
WLVxO1iMX25twc8NRkZCGCx1AaTD8zVJQUju/2xxtumJR7iSHDJVtVmsLdv9gWBNQX6LGEoEtc17
yimg2+ZYKJn03XOpXbgX4CFepj1NQmTDDciA7V7Yb4nBIOw35LzdsqbmLrxJP+P7Myxbr8ZtjJrg
Y9rTYaBTT4Ub7P76jELigKTIyyXSiXyymzkeeLa7Sn6Iq44hExwti728BOM4gT6ktR4KPH5DHOII
97WiUw3ea7KDkp1xLBAPB6EntRqpHIf12PiNDCiaJhDKgTQyD+btDqwWnIitBcb76RgiKR0fv/A0
bhQqN8y2vKbMzF2Ds72wBiWftfkBkmb4ochAnF69mcIo0JuE61cmWn9VzVxpeV0X22UbZ7Mrzg5F
0m2uqnsuSrL1/kNRcMZzmPmtQb1A4KfIu4b3fHwrEw3asRMjzaHeWeMqYuA6aXZSj+UGlvBKcsRO
SBBzP2cJs0iKsy3ckATKyq+0ESVuE/eejSs16iJJejCjVovXc9FDrsI33MkLNFLPf5N2ohnyrFF3
vNWsYGM5BJOTdiTuidqPnkReI5Zw8fZjuSfzNYLcfGeWPBkp2dMlSPUnuXGC32t+FmdrU/Pdj09v
8O7CzXACeFCBNryP+1HWxRSKdHVxJ0Rc6pW6I1Rbnil2XmcZBmumWREfOkWL//8aSHFN+Ee94wb9
kyZYCZ6gwfAjIYijW22Urs0kaZZlCueeHO4yv6roBXHvtmO/QKb8vTzucU5wsKW6ljiG7s6i1sTW
F7jLSpJw8FYwBAmV/t3tpxSlavXSLtvSJ2zVhGf0zuSirUwAyfHmUE3as4+Fa1N7z+1/XsgEprDf
msu/wwBBAfqvl/olXaeIR6/UfRNdfkxWHM1bqyxRzEdytLwR8UqK3AhR83VC/j64jaw1jfG9LPlM
6u7qbCwuw9hIJinXp0OIRdJWdZiJ+xkW+xY4xSf9/p/W2SrSY0scknN+lduwXIFIWOQR26LjdHM/
P1HbUDOJc9M8GEJnQ5UbokEKcpDo8OO0BArzJbrKX7yCzi8Sr3rKgmgBpnCqlqY3XELhOXUEmO1Y
K/rFJHpgfs5cIaFNBaPssVhCqggqoe3IcVmmirGknCMVsB8W11aQBfxafKOvhpPhKY8ZA72QLGwx
M9I2zmarDM8sCF3a6r7JALPy9ix5wkdMLaX1175V26KzBL223Ycp6vZIy6tZO+XbVkBFRZ9wfa7j
RzPnMnkYcfZ9cxqcq3WtGreXoYq9wxOSuEpk0T6ZuP/7qnIKAgUqlEY8fu5nNtMBdROlVqJ0z1o+
KHlCqCaiXldv3n5jhLYazS9rckXdrpIn7nQs5e/PQtK7HfZvj+v2S00H/CYn3PUFPe6rzt3XiOlG
LoDTzGQ9GH0+mazpbav5uIFjVvLFwWZucVQd5cUF5wBPPbp29m7ApIpwtUxnlPb0uZGvXaGJ8U7E
39ppOlM5XWutgPIS737WEYWw1mf9eFnbAD6v75aLH/B4aG+Hcu1Sr8aweFNO0CZAz+f5LU+YymUU
cdUCN2ODMJ36gWX/WLr7cH3llbbLNN/TVlMJdwHpBnjb5432zGPHMk/drV8FJnnwCFh0shJJBoGe
IeduF9bGVkgpucxpr39kvMu+vsKw776Lv8MUmmraPBZfDa8Iy6wewKLCdgRmcHOS3J9BJ4X4SkQY
MXp6SxSKBOrvWwd1qovGadplzax7P1konrS1r4W8HbCpMByx08RsP4c3SSqDyKRNoES1GZBF8ZjV
D7723SdDoxxBdQCXF0f+xJOdUoTcWCRgw2nC5Sx+PpjRerMhC4wpvKSERucD7FetvhRfZpoCZwkr
W8fqnKFCsjPmKtoWcVJCuXUW/rX2beYWj/RKV4dmSNoplnqWDtEiMKH7UuFxWqUcAcNNe9vo2NzK
W3viefeMgKOjSas+qWSkj9s5xdofPULfUB6B+bOqkMEQ6jqnKCytdk/7n9xGIZCo361/MeBuAvAp
uQVGhg+DZJU4uJkKw0G7+rAluMF/EUQTlDBpGwOOiaLuhWYc/Lq9jMJnRE4cIVUANpT157fzdWBB
toMNnFffEc3ncL8wr6Co88/8Md+BXL208nTy61mAACqYLBrel0ig3eoSRgU6c/jpam/xybP+7hXB
Aoo0xpVq/O+6xrqr1X3pdETklOpINeQxy4hOvkV/CL2YXG3RUv50tefSojP6g0pRJqCbHCEbGRfL
WhWDSh2PioGgJnc6lEatHg+p6Gc7pAbc+SdMsME45V5k9MWhezKyt89x+4of1YjMK1e5sVrBorV3
s2/QUioL6cfvGun/hZK/BBtNJ4iedQZZqfEJxHLn4OUOHk7MGDrrmr5+j/1xZ2D4i7Fs4zFZ77rL
3OxLaa/s8lhRK75Z+/CvzWs2YKlWP/2HpyGecmZ20ucs8625bu6vy1rd/8VUvhM2ecFR2rQyb/U0
6yXXfkArRxmAKwDGOOQbidmXv4F2G2renb13ijyx/DvuTPttRUPEra/7bQ9cEV51MoiAiOx89e4Q
buuOxQVnjVtoHOVL9gia+Q/mnD0FEtA/BSqy9fswoEuGLdR5D1lzvlR+k655xXOhP/TA2P5n8sZn
NY8ahd9+ysenTPnqfYp6hLLGqjAcKirQQF0lC7LzkgLSHpp2WwSQPhLC8dF8wiJtrK+Gn3kMKRer
/3NQhdc2IjAqs2PGu2+8ReOfe4p9ihPoiP/XCIscbogBP/vnB+keaaz7kAajnNsr4FoKbPzRx4kI
cfv3rzXlYVrl7eKDxARWhJfM1kxjsneFcRH5TIg7XUxUWcbkYbfM7LG9Mli6yg8YjFdaSd1Srq6o
l/icjGpBakcTggaRfjHKxzhrgxX31e1HMLbQbdG5nHE0PlKeVzYGBS2lkLYN88yA+HUKMNn89KLs
NINZSy2wICHrzlFQEyUdS6CNb4pYmyLg0yJvwWmUMaolO4nDwOHf8OLREcDreZaUq946cz2rl2zw
OCX0qg36dS6KkpP27ZYnnc+ZC5sAUB/HzNTUI+Vbx2IGTZwNCbxJSRR+Negf/H6EI8dLGJXaTs9p
2UKtrvpLEZya4LmcSDavaGkGGlyQLPpcWIsLnRsVck/x+dqpLW2QGMitkSaoEkZg2yLh9V1wYjlt
eSuScLBxLqOKWwnTdyaqxBzKnGfQO1yA+pRWUKg06o6m1HxXw5nqymrX/u2HsQ3hjVMSqTkz+yle
zVOtqXuZonB6eOAkFkpf1m7pnBTQkWnusPkSd1iIbxm1zXsfFqg+feHPIDGIoR+6A3jcmN4BqKrc
Hu2or8Nw/kkHJCxQDqo8Foav0k9Mk9SGgWb7l+TNZQzuSEmGRnE7616kaJmXIdyoUshqV1NRmf0/
j967UAIGJlU/W4QGoHmu0T5KkZRXvNxuJVxf+Cv5kZUr26G3bxVZmCod+NKNInIuWoRH17z78BgY
Y/fSxjpfO+DQqdRo1wgaObib69QQDYPouLEGEAl4XAe2BBeg78IchryagB68M5H6EUZwGnquBca+
6czU7CQtU+L/WfgSIpxFvbqAbIgTzx8x+HOd/zmWWGWWofH6QP2jLLaX4mX+qzz9n5qbiXbSgIhj
fkpX3HzcieE2TUzdpnCPt8TUHW/vIxBtC6PNnoTDYyRRxoZ/89ddXZnHBxXov/aeuFzVN+sQxrV5
eX5HkC2B8u+Pfe2hUbaC9TLVM4a60v5p148OIPAo7HxzaMkDNCjMiopBdMdqiXYHN+ZH99alC8f1
tPwOgOUJMts/3U6Ihs9cyNPn2QRSVBjCtHRXOSn2o6GbcBzQt0G8Ghjh7Ejhd5IL56fFMp17IrXp
yRAcGYPaIUFiGFvfm354oFKpcmSWSG9tB01Fx7EEF8FKcoAvkGyf9JXX2/l+SMxGFKC/jfHgrdo+
FDeMfyusJbD9M6cLdWBzcHfTS1Z8TakvVhCOmZyxnFfJh14zSohdcVPOL04h0BtxChJSl+HCHfXn
lA5RyZe8QKETi9ZGBuHU7dZn95fykE3hW/kuCrza4PLrSg7xTg29l0GOYZVjFLtw0KfiTFKpqBgm
sgD4TsH0Cc1z4Ja3s9UVIGH8T3nv7hIiRBdP2P8D66YU8wu+c8paUH4+U9Lv8TPysXKDrvyVjrKM
W/PSzdC1Jq+kwkrKrq2pEJiGjPifVLMP9K/EkjRWs8U45JsyZEj7dyhunmdmzu6nGUkH7pKLqsZD
AuW0jfay+syf5rfFW7Vr0G9SoXrMqWKl2P7J6zW0qLJTWZngIIpC+f6bNUK9cP9xmSGQszPzStBF
MAtmEDqqfSMAB8PEuHnkkxGA+YmO3hSslzstrZRRmenWqRoR9+C+mq4R21PJKPYzajLIMPahHY4I
CDLIO3ByjbmrI0qLbZY10Afgf6dVN3pVpGu9+mdePQ38PjuGcQdjGWPTOq/iCasrTJyGkAl+As/t
76MqGhNZp0NvhuceSmGycO16meEvhrvUeL+qYWQhSxVDpmndPqBvxL3HXxMheEvaJZJluAFUcRwq
r01V8yCaXSrbdPd/aw77LQOQnzQ8ldtSjAdYRDh78yNX3Lk97HLs5hzbi8/u+8kWuF19A0e4cman
9YZQbreKXDiAVhBDgh/fTvyWmiKxFBA0JsA65KztkPBycSOhenye0n+RCZjMeLHQB+7xlaHwKT2q
OGDdCJpe2PNc/TNkG6vlpcbmZTOHTtwlaBqZBkFXZYyzXPJMI3Gin0BCreb8G2r6UV9gEy6N9KhH
QbkJ+3ygTImWvIY5xtnK1ewefyLa/cyCSM1yVgAOYWoF8dHkmzymTTG6PfiP37UYQ5hEMjheCV99
nNbt9ZCmDtdqCSOvYCdlOKaGalf3aSmcFGc0COdouUjllk8++Nlq3xlByG31xtaOLAbZMG1O3Jn+
a4FnPHTt6JRK8Quuhoz9gZr5iRO23OuZ5T9dZ3ZaGsSOhPRadDgR308TJpZN0mZjvLJXstv8APF4
IkwegjAkd+WAU1AR4F7VSaktp2kdVgQD42HXH/im7Zx/Xma8lKdsbguYa+HlT4Z9Lv4ciYztFTp4
AlBgPpo5+Yz0Arytw8sdICq7iAjHzq0L7NbAvw1wharqiSYXAkj8stJ7KIiFj8w5yRVdUoaIYwEh
w+itFIedJzJ915690N/2t2DNsJijUgJT+ZwnZFNyHrFrHoJlvbC6OTL+Oz+e/CIs7VKzrIhDCFUy
i9Z8I+naT1PoDeaypc3dsOwWTT7A4nSDaiY3BiXPUEoYF16OnVOtbIlGWBCSTEcJoi3fUBw8W1KG
ie8Saib1a9rKEOTiiSl9H7jm8WpfoAR05bO4X25TORSy81NmQL3gbV2583rY+A4VAi1rbRVuf8Aa
kxu1fLII8CDQvCHOQi3QXg+kSuF6jv+Pf2T2mJ4Y5n5denVleR+2K3ezSUPqKzXYsBNxKFQ4Et/0
5aLvhkeCcxzm7TmR6wnbx0JT+huuqb7aur/qDRpBctvNJsMRUX8SlwNRTbm86fHeBilddNm2Tu8J
bBFEKnzTXScXHYGCWSVeUnjTMT2SgQoXZuOodL4gyb5uYBtOwkTXXaNHYH/2jHM5BZNWdspQAiQR
wWDc3O+Rw3pTSV+AguQLhK+H9EzPOSElZE7bSTlqRqLRiWObvB2Z3jcAptwKxn7GdKU1GSg8EPFd
6IkSjautHvLtwbkg/eQXDf2G59ZI3fEnNvOlVJsQfqS49S6RZ6VkEGL1AmlE92EBhjTRccN7VcIE
65092n4pGJ5p5bscZ2B5AWut91yaMlVWC7Or89jZp5obQamSA1CD/0EqUGxFKGplsiEBBvLpZWb8
8WVthcPBi40MzFfqxB10hx+X4KSqCACZGPhbqwAL/FBPnmpnH+KxLKrE7JZAYlyCdhNHpZW5Af3C
jHhHEYQHEZtGWDN7a76/AnPuzsNFKVjBMCdeS6uxC6fZ29TEgnFLlhkFVx7kZzQcpM0xanGvuDzP
FXVvleAza++bx0S+a/z5ugYaqlOMxklU1ajvSlN7aKwybpEfMCV+nn5waaJdCYNTV2ZSWNqwY4XU
HfvE2Ta1DxaYCoF3cAbUkQEzjsTvFyon7K+79muDQlfNTc9m/EhE06/isImuzz+ZoAMXzSB/+BY5
8jRzdF3TBcPUXCj72FvTsKNRuM1bjvJhzYdc6RqFsdJ4wY40gJ+ZRwpqykfx3GnjPL+KSNWs0Pm7
DUjHTNNACB1oODtZ3kP2anK7j/1NR7qVTXERkOW9YXpMVgsh430CaRF17VxWVZBJmhUMRXaszA69
u5NzEzE+CZpGX4/lntOJshEirquLyVoAwSY1w+YiF5R7TIWFduR5+HprE6afHTGzcyUHeLViBmLk
ZFAUMyToSe3yxTBU0gL4nl90xwl5JluC/ywkbT4QOgeSdGE6Gsy6hyIZpzRwrofEUHjRnsR9qxNV
aOEQxRhijQ3xsuxhdmV78VrNMkXog8ij9KFdyNyDia9JJN+okGwobEa+BXaE8DJHJZMpigb+/a9x
2i7LF5NWGqBGuPw+mt6aCJiBBYJbsznC02a7usiM3w0gx5VPxumF0+2JziFnMY0NcQV2oMX9+Vhk
bntPMrHjj/qLvEENktGbl6yG5jidui7bCz6quZZib3pG72BlrU+R19XwbgFx+0fwFn6/UEDY/2Ae
nyIY1ukJHQmig7DZ0Th+XEYxQoa9g2XgT7i3JU8eQ+dfOC5qnO7yIujMFeFAHgfamBIbF+UkF3lX
musjCEhKHvLE22LLufCpHAalEK2UFnZCiHFfFZnzje0BMiMpMvPHWtWCEGGslp0zkuCYTjkj8NJ2
Sq9/oYxOjYez4ut5GDVpuBLCqgoL2xACZ+2xb+LCIA36w2+fj5JHgz0QytM4cn/mFsxbnVdsR9u4
NlafYEAJayudMccb673KJeWa9Fkp7TDwyewxW7Ng+9ZB1fSwMc5tG3wCE51PZQ0g8FGB5/XJ1x7a
23az05MnX4Jt4JxLv1mQeIUfXlUJ5UsP+YYEsNx+EHgeyxKnZq1+8r862Qyabc/YOCqiM6nVTL9M
pFHR44YAcif7V77tuHBXMEy0HmNIlD7FB5E1KepOUwy3KKXIccb12OBWYKHGiJkTuVynfu9U8diR
s+RPhb3xq40F7Ua/1CLqmKvhtoX0TE41ipguKs/VP8kkydfST8+yghAWvslwkzuAy9oQFK/Am/O2
cVIA7DIl/VbPV1qesg==
`protect end_protected
