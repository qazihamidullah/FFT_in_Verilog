-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
i87P/yv9D+pH2Uu5srQ2uKkgrnhxNr2JeV+ygbljPW0qw8H5G891jc5ic7H6Nddi8hFXauJpVHNF
Ka/zpu0yh+1UbeKC0OdonpEOlF4/td6spfHwBQsBtYLyD26aX+DZnn4jHPMHybDdTCRBy35LllEw
wcTLuPGouvf/d87lxyug6SU1oV9w4DNHhN8STxnPGL566wbU3WQ1nwKJm9i2ST24Fu0xAaJP0B9S
G7wReTAZDcX5G9qZL3MlMo79PO334w1tiq+j/QZtGu8hqFZZFI4YopFUjshWM6qx9O8DjoZhJXFc
RxnzbkQamPLjPSlrPw51XlnG8TvfuQGpiR/IZg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3328)
`protect data_block
FODzX060qn/hr0iH1WI0telMHDENlsEHGV1SgFOaUH/W+weamT4S2/yPbLw65WF82hTOhNkUwomv
AosRC+AU+6jAjlQyowRsnPPOOJ+h7h0WpA9rmdJUpHHJd7MdMVjjwcwsfx5+ynLu2I0Qei2L7wl8
gfGGJjXCABv9nvOXNZcy5LYDFNGhTgay1INHyiG4dLCUauV2oTRYZPjLJvpoSHfXsxP+cz1k0yhB
E+wyyk5X8Dt8AAifXLdpm0P8nxMUCJTj/+uVwBRY+Ra0fjE9+EvF0KMFtxL9JwBVEBJLgB6azZfC
ZpvRBUkQdivoMOzO5mD22+19nxRmhwZCsVS0juTyAIWs8xmWbM7qTChxp4OB7kW0Kf1cijkcRX9H
X+GGfNcNI25hMrYMgevphYtC2l++DYSEZTnpwSkWPF+KcOl99tz07O1pxg+FXu+HG04a1+81ZuYc
i2ZHQ3kS8CoNir0pMqUDWRqjsV3JUCqE8XCIaYTuF8YgGxUU9h3mAN1XybCzCkf/NIOClPkGGQse
RUDFbX7Xq6aCDN1xh1QEx4OMPOC85Sa7P3j3F2S3XrwwkZjiJm+8tla/Of5QJa/ngH4xBWqZzqxP
f/YPnZzaA97GWH9XGxUX+nENuhaRSB8xZqIaCrHcyk+Vwdda7pxZJbU3L7yNPJFkLFMgL/75ttPW
ylif5NrPpLuo3wnK8y/sFwP2IbKQlugyGpSbASYE739xQ4AAWvST7oY9P5bInnagNku9gCpQNIPw
TNuKyrd/faLund5eqnUgmfEKRYLDgL0Wpkwl303Wfp6sConMCFmRqcuCKr/WWXBDQi1spyK1HcCf
+YLbXHiqQ04PDvqxRl9Ecqz/HKTrYCYeMMSO9YjkrjvM7s/JseK//RPQbm+xROUkWvjMm/0zg7pz
p9/YK5JZVfkWH+oUiQu6lgl9f5Gc+mransLCHY/lqJYc81tXMMtl1HGhBunW08CsDayDMiam2GQ6
hpIYkAS2V1jtbf3KThBP2UsnKSKOUk0o6vCn9bnf7gXiVOqzsL5jMAEyVs6QxVY8tTwzKkZZYnfU
fBnl5VlQAgqqcLv4v1MK7hQidtyTQYkzs4S/c5QJsJIVW6vpU4+wfbksbGc0WaLP74yJH81TD87U
1U6ukUGY17tVtggF+qIjCW5ZHg+TFuw2yhC+0zcUvXGH4NJJUHxd4GFGktFOV9rbJcnkZ4rT/Hx3
haFk0OtRqqp2wbfKBnYsM3+GTcfXrKZ5jEeZIH2Ik5Dne+5bSAxmNwddkuEzPqr4y1yW4Tkyz7m6
xo41wOiFs8PxYjVtozBoOrlvdtxk8k4NNiH3LjUKECt1tTYAkO5wmIe00xqGq6gvWIVrPMYEH6jx
ZIi0rqlYchZJPRDJFESIMCX0fYSveqOBDls7NYvYJvqF6Q8PRkhUQprfoOpLrLcsNZ5tbEncA4du
p8yC94jqg7S24fg//Y1NI9+zAiKOS4waQuUzzmuNrXviebCMQjcDi5DewaDq6ceYcZJZC4yzYnSE
lQtQoP36BRdGrUtlAD0ajY91yBjfX9+VI0GJTtyPuXhyttUwz2G3mDGL/sE9fZC1IHPDsovdCAkR
ZO6yR5HTA+X+y6eFbzhaRTFw1TM/J2B7FxVcqc0axmOEch5NauMdABqTnxx83hnwlA0Ab3IY3U93
u+nv/Y4WENL337MqHbLllB9jOIDnWTC2X9DG/lLR+HzzmsoR0l0Cuyz9gGwwEQdVXgEOZXC6n4+q
qohBJCEzXri7S0rw9WPNIMO2CUJ/Au3+J+DUwgtJ2VU7TePsBz5w5/2sK9IvTVqsJvo/A5QeWZOY
KcbW17wdH958cqUHsz3ydWhBRxgZ7oVzRxWbwYeJb2I7OLwsxx3WCS9cnXhuICUEKHgFk+ZFqTDd
ktvbfXXLhcYHpawgOY8jo3QksUUXmMuA7ZLJDXUlvjr/rNjyJNLqGao/MHLJnZ0Kk07oVOdT4Od6
hqPEK6WanIk2aUlknpyK9YFg2e3wd49icrEGUEukmK9mL6jbUzWq57uJzDi/G9ibsbcO0qsYwpQ7
pvwD7HWe/GIDRECS4sUHRlZ3maLjoDbAiUchN03lTrw00YJRPhfiAazuZjMdC4k10PTWYoN1fQx/
9U3nLPbWkWIIzbq5IvFIK5uaI2I4CE6MY7U2islaQaYzgfkuXoY6I+z9I3Xrbo8qPWgH1Muyil7T
vEhyO5MzvPR6FK7sqYU8CBSC+UKMMiSTSixLuLmtW3FEe6u0Z7ELuawsGlWPIkSIyYgxKjgjMaYr
yQwHyEhGqC+7hm8Hnw+srindax3vkpGCjcCHKof+T6oODwgB3q+j2NrzLNhQKhBNoNkOhvOg82Po
YQVFos6Wxbuh1OzKOUp5ZrYdP0+bKxbAtGCsCpioHpM239voFQhSdIjIHJ3EUX+Rh+2MGUSS36nq
HKgfbFE3UeBX84ThonuF9fXf+3z3Lj6PbvcjFyIg3vdhXKZY8d7FWfbztmpU8oeApLe131RzMWpA
sTKu83EdmYWCW8qMAH9nDD0hgAfF37g0MmtkEL2r59wOCmznmS64xEUqSknnAd5D3EcP0uAZzh9U
vDH61Ap/DJJ3ihPWt3oLG9M7ZFdjqfwG2u+IYiCocYo1buJjTt1wsxyqYryiq5+vBN+2wv7oeOy8
3rPOTOxE4e6yx+IbhsngC9jTL8/jVNSnZO3KnoRFBEJwOK43mWysIdkrTZlWUjbjYSCGFoYmsPag
UOw+wk9W7ws8tCJkezbk3viWizvx6zgG4dog0FXb6qdypGG5erw5YPXJW7+MBZFNFl8uB4e8uEcn
2/QEY/aGeK88GGEh12ap+fF65BT9brwY+f5yFyJ5vhRRkGsVPTKlAeVdEwSu1cA0W4w42DbE6meS
+KH+DAPVcRRCx57mgGYnvp0Ct/b5Y9zKGVGt/JxVXM3DZzsonNSjc2IDYUTzs047V61TIJuM2IoL
J23drT0QXBOcaEiEhkmBiTblVyhpDS/9SyAATuzWdfk99Z9R/7or1f4cFBuzenvtsw7o2Z/1oj9V
0NPYML7MS2phUIkFj6n2j9vZ0irDxcw3BW/wvNl9fKgUshM4sFUR+dte21hgmCyBhTzFpNd+dGYd
lRqxipucCaUE4wDz0xPDt36WPltACpO/hinMUlTAMdRoHQC2/RAHE3eH08CENK5EF1C6olcXyYPO
+4nreoGFrw164Brdih4OwB7gHRshKskYz3juOJtSOhBbvMqvuSKpq6uK2ubRBWGHiXUHBj4SPMsD
A5Q8esd2EO+UkhUhKyszdKAC/s6ZvRVMP4WPO8DIBsJAuGho2ZpoWyjViw/Nw2QFON1JW0Qfd3HR
RFEAGTV5zVv2hhqV5QWellQ6h2C6xEG3yw1bxIm2ubhNtyXgJdjd7oPwKzS/RvjVlXtXJSYnxDu6
Xwev2pK+UtpGyZ5sNK7Tk+pSHWNbvgKAcO16AQogmyupGMKhjZWoCp+kABh86pqMA1bPiWDWbFlu
CrYt6Aa0xgQNJy9HN4fqx8NkcV1l8paIOOUo9T/raJo9O9X4U/cTrhJ2VwSFJlWQ1eDFqJVtkj29
TA+d12rRrpgO6ZJX0T+ibuwcoYNmD4fU1frqC7AzQEwqyEGHLB4JUq3AhFU+gDKqXJbyB7EEBRb/
p20n+WS/7PjbXkn/KFNgHOOVR7n2u23uioeAmLeDLI3LCVHWCH8lfKOktWYLmev6Z+DlNVr2FbqX
mdtF9qGLDrmxrgvcOC/mhqFZhx1rfD1bDaCbvboRp0waIGjRTcsaL4ggncBnMu9J/VzGiSE+TkUk
qzUbuS4bcO6hDfeBnm5lO0e4xj3BD4AkwSH7g02gDZsLKrcIPukyH2ZjpaNnYjMRe30bZ7ecMLfk
X3iGTpSs5sHk8OiGHA5XFXHp/ZhptK2B3qHl5iAhBXud+de8WLIuMhz4SjHXghews7mdA/myU3G5
BAtCcgS3vrU5MnFt2Z8jGVoGx7Nup6A3VHWW0d8xUDP27ZC7uachiEfPKgjmyEaTsb/TbcvO4se3
UOV0AwJ53lf4Hn7HzpokG7TtebV1q1sOhmtQDRMHrj3CtBVMNmmd+oc3aitXDW+7eEjOdkmyu5n8
zOsH2ILkvkMaAuGSOv+ZmA8OWYndYVuNpI+LZQNUwQMEFg9fEkoKK0t8MP2yzB0ZrJFfqNO+iIzz
hFKIxl90bbl1zdRNMmDIKJuwx7YJynwETPAsjQ1S2NOVreQ8CsafQt3bjs9aBDtqJ+Kq4CWcR7Rd
6sWCj9Pz9Sb+xdwzkWhG4/hIyMKzvFh/FB5ndcTF9NMY1A+jID8LBMJwSS4kZWqAxfmvJeNDrMva
pdAbFVS+f0/NKUAfVhLu/AJmTIRfVZbRQrV91zKUMmwrA6jM3P5FtVKkF2+y8gM6lsAkJw4AerEn
puIS/qLb3tqPz4NIr6En8+ZxQScudA==
`protect end_protected
