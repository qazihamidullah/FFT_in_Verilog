-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UZ84mbd2gObiHNahuOFo5sgcMg48+8JL7ObNhF+8QKSrFHd1vGtY48aZWt7ex0hMC+vWAXKEGnuW
bsQGICCdPOTKkywClaK55DZSuRWS0q15y5nAXJKbyNIB53A1FT7o1RXPsAsHeOCquJBPsoc/Cb6F
PIyN4FRQ0xV/u2WulT96Qfv1ZRdQrK9FUNNk5S3JBUYo3KboFJgFl6m9hfky3WfjQvbJUa/+fgjm
7ftccIZtdPfU5hGjzZ6SdxQBv+LiDvYnaAxvaSbmgedn2MeFS8qqDfuT7mW5Pc1LnnKzCF0v2RPj
XrMJ8hZCs7qyb6OEzV6pmDF9lk6byYnb/wwW1A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35616)
`protect data_block
f5Uh93sUH7ne14KIYlKzRFCkqyXzu20c4b+EiAs+OQ9FooMkieTQs0Wc+0OG8Fd9HoVu3XZE2bb3
PIIn9SIGRaAX7XPNlxTcVfd7NreAZpAlXO6a6Xxjc5sy7Cm1j5/t6jEo4VVAc5ekDUeiuilCRMr1
JhBKnqIrXBTkI/eCvMG9UXiWBRsjkOV5GGqB2pq4sJoTlshzuGGh8r1C6S+ZYXA12+AZMBSofses
dm6pG39TYT5eKnASev+Bkjm2ZxZmTty2zQlW4T7PxJXpnTTJxicsghJeS/rWuwM8I3AHzJ5oQdda
oYFYrWR1obhfopcJyTQvVFNJK8c+KFLfFR57uh2w2Tz8ZxD34nBe5fUbd12KTD0JmOsspbCH9Kqi
18QXLmPuRwr/0jmhlEZ27IPoWtuxpEVvhNutErfVAKl1Z2RdVuyYjJF73Otflfeg1Ztppg4oyXOS
L7qO+2BmQbKMfR//vatFNynr2wv45WaQ5xw1R42Lp6/lDUp631aiwa3aChDXWD5uBN1inHR22koH
PKxLX1kAn7YRsSgKCh4CFQe9TTcOe2I+Cmw32aLWCwG9qU3WpNSLU52pJmoYdHcr6ZsoKXYrtkq/
w84UWXHvPHasrI1LxIoc29sv/1OA96k9cW+jYdI4b5B/3pDa0i0a5n3RWbN03eg5rPRwg2z4llZP
aZm26fz/U/WLPdxjjQ10/0yeNPiBXrf3A2re8RiP2RA5jXRkkXZyQ7odPdQJ1FSJ3SdoKDXD6q7m
OEHMVm1go+1Lw53oLbRiOaiBtdVCTnQ8jQjMesDIl0vYouwmU+040BFqh26nBEyTWecFbrfhMb15
U1yZ9JkePWEFlIR8igPZDfqAr5eXtwqzt/ji6vbOUSVaAp3IAGMAvnmmKhuYQD6giIlvua4wd2cU
xxdIR2N2tDHcxEXtctl9kz2IlyVyGoHINhefUZRWTJWYt2xtwq/UYK2a6tXjgEhca3YCbi/WsXjv
riGdj5RZOx8xJFOzwwug68cjlLRfKa+sFzR7Qd5CP3RdtqVCrClZ0Nsom4eQGUUoPJWg+FIXf8jG
9A/g69Edz31Er6JWhHfylsno+L1NrOAH2K6mvh48u9l0Ez1DHxMKTMxSH6lFdprIOIMSYfKFsgV1
Hj6gQVH7mvrIlHxMfcwb/GJeDs0i+F3yiVy9lgm+/kjaACSVmsNKg7cnM7CGQ3v38js+s+5c4glb
i26mPyzSuOEACTmZeKOhtGn/Ll6e3UVv8/Me8anQqCdkrelnUXF7Ctuje9b1smJHtZOhD/1Fz0iE
N+HhonC9Xe28gjKA2KfIysCay2rt82eG02+zfKYV/w1LxD8tutXuLqsxizSCBFMI5zfoS8clIzhy
1JB5zFoXLVlV9sKhvTfPcXES0yZ9NoifwQaRoIiSEuqcb/FWkxVkAuVu7Kd2cZfGMVlj7fu/9G3b
/33hj59TS+m2kTpl43eZFjIiUmGNCET5Qsc9VoTisuYNccFy0g93OktF/nntm/1xTVgk07l81J8l
JoJgPwrxwylBOpKuwqB/DcmjEADxAVDPCyBZ5N7eqja8TONRxYb3biAzv2UzlCgqvcObth7T4NaV
0pBIc8c2JKoM7wSa1X613Q10dHjDjrnRQbXZXqTwnpYyUfwmHQibBUMYHiDs8XN9ayRhAbECCT1y
FjiUEKymDhmG+bTZHD7OQmQL/2LCpcnkP2nTgiBEFoDiAhfXjzY2rhjJdP9ywUrJQIJvikWFTtXS
5knShXt5IysToDb1UgbwPeppbxJgH+TFGfYk9bmIjpVrbIjooF7XYeDPKnZP9OBZzMB//K1oXXv/
xz9uhiRg5xSaSB7wBo61UvEWaqBmi+qcJwQ2Pmhv9yPCaZ5MuLyVhYHxt0QZPVd4Bml/t8KihqzR
rA/6okfweIh+2WamJOfB/dOTtZemLjQYHpFpvufbOIAUx3DaeEYqh+o7Ya3fNk734k7ALbjxhjxm
QTpV+MJFfZKCwzxPGS0ftNyvAIZEgOXsMrtBF+tmNs7zwjQDvQsj1I1qUNm6t7KGvC8isfkJ9uz3
r0IigIswB0wxfwDvRA3ZU4yOSc+8ehg6IabrBg3wCUN51GmJnk5T8vX1qUz6xzNVVbyJcCQy7Yl4
rbqhPpM64pZuAl9xgSDgpsKrX8TOxIB9oQBif/jGQLxt6H9xswwDbNOXPWmH5Szp0s6akmCdcJc5
GblwhK7L2BzXOgY2tC2JBqu2wwkqQzq8rBLd7YWsm4qWovecVP7BqBV5E7MBF9TtVVO3fkWRBAUU
m6tbnET9pjU6YGppEV3fVenZG6ti2pPUI38kGO0WX2smZXFvpa8EKmC5v1hqkPb7yZZ/3MobWx5z
vlIyoN9YK+IOLZaTJNN7sCKK8PBKCR7CeasS7jydGcWrn597I7mSDXfnkzCQNlk0E701X1VLlJaz
HlsghE1cvF3+KPfa38GLvIZUl5IsHZG5XOMevWzI12ICs4M+kGwjkYEh09dzBprOtCM03Ll3Vsjz
p+PdwlUYNi4wjg/Rd3FGbtkmpEwJzF3OM/+0GLYj3y/jV9i7fcmHvFMDUIh2EiNqNdVeOmc3llob
3JmyaGZnKMrHy9FTdsdSfDKQf9dhN313Mnr/1r9mkZqb5h3A0eOYdpPwNdIZxSa9V1cyUayDUnla
dcgdGvm4rWauKblcD9eirXobLst7tJbJ+rd+D5Ue8p0l0RXKbVNQHpnH53RVLt1zJkyAlV4dWGEq
KXTw3HK7NZoL3Tm1dP5QEMx4DctwRroThxVyN4yxi2YJjPcS+mNPibCNx0OIUSUWyxurK8G+zDQ8
i8QH+z8hVVivvXv7hSe7KGA3Oblgqi9MbHtV8ynleOCRa6M0TiLSRrZ8KAQxeCnY+xnYZSrm8iHm
ScaPLhhmfVSzr+RcySJcWsG/GcS6c1VNY5AgFWyNbyAki8vRpo8ul4iH9CptABlF7rIhr7y4SBhB
PkYciLxGX7Ba/cP+HzLTOlAliClAB3/r1FQ12mjObRsPil9a4SCzfdVWyZvPdeviuWydiJyKEP4p
REWmJp6FbuS7YMsWXLwDLHC2y00gF8pHy1PwarH7dQcwEzHizfACkdTEuBoKApj2SdECAgm0pKsq
MAaP0JalcB1t2XrjU/75IV1cLGkigHgi5qsqL3fVMS4M1j1tlkb9/wZ+mAZJUeKR6xc+otjlcNvo
gNJo1qs4kQ/BOe+6h7dedIxdhf59BP+Yf6D26TmzpgT0opO6ij5d6RkwVAaVlw+xda5dTiWhcxq8
SvvCqM+phll/PL2HVu+8ga50r6XklK1xBKmHiL+9YxNoaOTX2u03BJb9eYhV6s95qsFbAkJR3Cj6
gEgqkO4EsDGVlsZ8OfAMqJeDCH7fodoBrBHBnEEzFfHwHbBoq4HlvVd1ljmf0FdG1tfcUps0uB0h
eo6B027yxCbkPc8tXz+S754iSHYyySOI4+fr4B++M2KKFRJ8HNSXCR4tXNq0RU6cvH3jXfNk19UJ
ptFTihY5+98WIayVUTDnSGV+dz1ZMls5qMQkY8D4u4/Pw3YgDDC2ABVA/YqrpR8zHRy49tO/b7xy
yRKhrZbwZBiQ2FQKcKn87x1jV3Re3Ydh0zbyFRnM59mr1yqHeW0aeFevFHvIrtxZ8ksayxWaq2vL
iw0dlBva5TdXRh3N3kV5R14190GZa3qtFOL+sdyjCKsyKOEXlu9vaxdY4/HUGprNJLT2tnQDU6sw
PcdiMtR85Qhd4KHZRkbXVZp8T3TAgdyTvgDRgtKXpBzXbgP9k76bwEb6h/5NCJemByJs21uGQwmy
bOXrwD+h1xaKDTGRGnHuMU3gy7WOoctL/dlmxBc/Jkd5p4db+jfmJmxJNMycp+tCo3lK9wMbzsd4
cTF21u048oUnSzAkBp8xMJVYm3bzGMUtWPvfRUbDYi2NJs0lPIYIWD21bwtCczPKzFfwRIPDy1IR
3Z0b5Kp3xUPAcEiE1EeWVNkZtImIJ6xWNNopiE89ybUawa0cX/F6qJTiKDSFcf0akMkGkb8hOWcF
BnKtsJLbTHDver0m9+pecEuUNd2hJL2FRhj1LCztXqG9uEI+2RPe2Puw9v0I0IRpM9DW531qmwQu
Jip6oWL8+Xz0X68H3JgZIzwRTkFvHvHP3Urw4A3mjno+PKKDwxToYLkitaGC+dfYRFx4N2eU7pl1
QuLiKWf/nTICBA9pmHD0U2fJbBJX+z/4fJlevjeMflRxrOmTpiVQ5igjrwDIdHtJbBbQ61V/MnSJ
cVUynwHDwKzh7Ik0KtzVI0StasEOj1bYuRsM9n5aHoEVCD9u5LqGivn5/CmIuG4gdSeMed/uQFZQ
czf/avJ/XlctluPk/V6ZRP5qyGxYmk0qkZBAmA/Q+XUduVOO+0pDZPXqJHktUVCeotQcXWamZsXw
XtONDN5os+E1eHxjIhaCh7apOzzQqT8nCvVam4Xr+WIGmGqGYMz+20GwUe4SYTKW+aVIjHfCiifB
Vi/vnNCdznUvj38aUJxItvmk8lcQYwpkP4CnRq5jAN+W8wHzfbKIq1rp39B08yjagair0Qzxk/f9
G50GCTYdv4f2x/3GGakSH3iSFIESUrlYEhPLTlTccxcGwH6sYHn8urawVyvSLEhIflxEdTos7sTi
lHjTvC/JbPIYSuKAyDjc6iSqhJpKvgAw+RB9Xf1BFS8CO/xBuaqmyeprZzyRKGcQjXArNSYQiVNA
UVxYC/3sEr3i6nA19bgdo/BLo3vA6/NnBD1ZfPcDKWs/muXCVUwdwXJcm06bU/3gx5pW7qoMNdV1
V+2LlrjELoMxuH5NcCZrirlM7PCglkKraye9zWetq3EYjcfzl84zcYjHgbm9d3NrDqMzT/y3M6CJ
EWKCXERxrP7JsE9j2dzt+Rtg3IF88ajNUyUW7DAv+7iRGIkevfpQ6kBAvBtfxZ8w3BZDAWDbMvxG
Ulx0j5Jv60vAG8CJjyVWTXaOXXpIKmP64skzETA9qUGyRBD4I4peQCaCrAPYT96pzK62p0uQqNhD
0sFShvOPlstnUej274eqQeLQhbHRvbslFSZORidw6eCBFVIGZt5YfNCpyYl5uZHbLc5UgYYo1wk6
0dC4dW7d5zvskwZqsryEkWqN2WhANi8Nm+mSOf+ZyT9SaN//wf+s/tUggx3uIv9FEzUKqgHIugcv
LibeT2d3aY350/ywNxa62rn3MCM5gdCw8Y93T7721qdwuH6CrFWJDf7Xom5qeSlQo1jIqY9OvtrA
6YWIPZwGZ9NlNIMscD80DoXef/PDkRrH6VGqckgywJQRN74qRKUUgoz7zxWb1J3L6l/UGlFVOnNU
HwG7S2LX8eTWJqhUIccB4JvHwV6E7aCjOYtJuybm4SjdgQDQTrf6/737Ib6RK472SNIPBfcW3Jm5
LSUNlS79K3/AVnkw21A5sEqQiqiAPhOHifuIp9p//15fcq7LTnqdySs9b/hLC0On+mDACSn13hje
ipWpd8CnwGJIZeZediHFxoJ+7s4AqBzUvGtS7gEt57LeqFRWOb4DtNYECwnZ7tEcNvxF431NypMP
HdMAW4SebDMMqZOtc+CRdYSRfVICoPAP0e4AlbikC4fuf566IK7+A34qKvfN0siWPn15/MWFjHly
QK7aB1u/2oON2H2FK61hhh9ABM0hW/TIbBD6Yynp9etFj/4aZW9HXZTT5XGCDEJvZWx6ITtoeD1Y
It4eu0WykKdkoEhoJvqCc+BPdnrjpaSPT4IkN718HlsR4zm5dOJIqY0qR3/IC1Ul1oI35taOsSxk
u97npNNBQ65WB01sTcx8BDAERAlHOGGuIcXiFxjktMDmitZWlE35muN4LKkvKSlGAAANTQiZ0+ul
+BlQdpYavRVuF4YfKJ+MfOf2gByZZXkRR422rvSip8msQAvxbo2MVUH+xuz1evTOCWN8e59LzVRX
0Mrogg5qohAVHTiB5qC1wSErgP1dj6Zi4llIFqkN6zokKbTF1bx0oPRneIVgdKFx+wFo1i2ZVdc6
N8+2pUkVyOvwqtNhOAs8eYmpDYbJk+be4muc7t+69bwqPP9RQPWfLLz/cTcTyGInKL+Zd7eJIZ8Q
e0g9KqWKwXYkdGZxq0vMViRF8rYkhgEkeoq5NpoQsv95EIepFBGoVkmfr1iHt0hRqCeAINfcotMl
KWprKyPy2sAqeHljCPwfwRtgNBeCxRBDGS04+VROShS9MNKrpk3BIt96w1PN7bcaS634hc8N0i/c
Rlxc+bdn0D8KWOK6eO5RqLHz96L32nv9Liq0IErEhyzta3gf3YJmjYGXQdFCsT58fuUmla++PhR1
ffcax1QxNwku+fqb1pjjjg/gmgO1P1xH6P0hDGJHGch2gwIUutkk+L2p87oYzH6x09v7UHWang9e
J+Rj5P8Zpi1Ga0erX29T+6M4FjVYA8tt1nIa7S1sX+JDN1Lc5O59S9WPt0Q3MdZaDq6fXi9IJFsa
Hb/6v3jILrwOTRMGmZ4tDr5G1to+n9i7BjmqUrFTAsEURlewvx07/3d1D6QgYDmbRamDVbQFHxaj
af700PyQue4KSaQg4imhLLXKe0XSrwPDfjSVCCurliAv2jWaZ6YwKjTrVWgeyRycbGWZbJVmxOeo
CBiC/Cx4Qp5Px3NS9QUDJWhvu2gD0tXg+hjv+7MuHhdcN21B8fnYGVkXoJkoOFg0R8H0l67gmxN2
6sjKDZJ0nONlRcfXSVxP7/uCzWjWOwoX8hEtLzlXfrrQCEsy41tljEs0jDhU48vLc152lXSfrj3U
PAxXvSP7HDjoqC3d5JRBAZVDQ6tHq618csTYWylCrIj6hx/K3oT/9TF1j8Ok6u2AH+fs+VFF7bLK
Mn3TK2zFWU0kpMF5k+4xG27aiO80bVDoLXr7y5JBcaWTJhsyLS1TXEN2BiZQ3NKnbcd1ofLQQJmi
zMehad87H1Tun6Qb3Gz0KMrOsydnGO+/CWwxxHlOkM05m1pC9RJe5fs67spd8Aqph8P51J0KnFO7
UvElhA/D+MzMLuzA0deKe6v1qSwl7d+Ruj3MP4cmztU/vMu2mh5sDiq+v2Nd8T1Wi0+OScVlvA3a
Swt/P7fkKHhSQM2uaZwt5uxxlCCTq30VWGpRoAdyGorWwkUtJcaULAUyjaJOGPjSbuMOzKr2ekBU
trM3hQXSrTzC/VE4H6XYAz+kVpTwvgCVVq0zxubqSpkhMIp+H3uF4XhodRnX4AY6yFmBigdPrmCv
5rdh5PeOGn0w09L0nPvStvugaE2kDViorqlyPluX1uljOraNiAkgGok1End66XF10s5IxsspjYSz
nS/e5wYUUKecoD4w8CmT16okkmUH6mHoQzuo4XShHA5pjnqIPMn6agSOAY4TEiy5iNlpf8C24B1j
IkRsZu5wI4GpuAE6QbENhmdiOqmgenRNkBA6ijsMR1drc6B6/u4LqRdz3vtLdFnFBlUPlUsM8jXL
L2pl7POpoXU5/5P29nOC6h4UTW2548PiI+/g8iqhIZTohGzoUrrZ52lf3pH0PfTLde5lebo8G+3M
VMkBRbvoa57hyORXIKs6KcwBYo+cNTVto1XuHRz86o9K7HZqZwqnaiCTkKh4u69HJgL4PV+1s5w1
FFYIRltkxbC8UYU4UNDb74uYBQF1T2NCVj0B4gyb4Pk9cFzkRsOxvo1iKFBBR+cE5gvwEVHNndzP
CUM6KV8IbJYgOby3A1DIEm2Yag/VbeW1qAcppkkyN8NkL98AxUwrDFazZjLCHkvHqy2K1eCJ5D0g
VNLo0K65XJpM6NIoO2l0PIoWWOSSxTRzK3m97eZbOxUORvM0FyBAOu85CGHQOvNTFlj50KzNd0HR
mXHGzhbiR10gyx8Qcv1PMlwB5xL12juC/x9UzgMIYLNE0zXhF4JpzY1jAasFnbKg6nzRoAbeSpBw
fts2ijnjVwARHfhgk+uthWPXgp7aAZ1O56wrZip8JsrFic+MOsqniF0D4nfqFUglkdGK3awtz+zk
QTKnvgwZ5z3Y+ff9W5sjy7S1aj0y0RZntwh1lkkmXqJLp0E8SfY0Tr4eKwGAn5dTaOUGM1S6nq/R
PexdH/FqcYPeeXmcHHJ/83xYeX92x2Di8YWRV6cAruMihSvCpLTINhhvG+jR6FpqqrLa/cuaJQLD
KeSOWQOnOMeSrz3qnIDmdHSvYMWqvWUoxaVDtdvNNlujwCewTE4NGmxyiukvY24ANbY1tSd1lp5C
Bw8sT+69Ipji0X2bDauNEbY/HCM7cCQ9vdRJ5pHN5fduQD3JqVuhT5q99I6rdZrB7WjwPVoyAtwm
13+doCGkcW8Ku+bBxNwYdmryF2iZmjH7fthLMRcENPD+6vJwSFf4fKmdUwr5bSUzkkDuG7lJyDdx
xMvOdh09+gd+/ioPFfVFzaAer+U630NyegM0EfHVXwX7Cf/AhmASx0eFpcL3FKQaMbXjGldJ9Nca
FBc8mf4Qzi9+RIH1K3QIIM+CbYfwWlS2t0QBgtou8stH9OORg49PJ7okvNsfM9bxaL3HT2HpRtfB
HENDpTkESdt1NgCYon2G6quoueFTnH06aZcMT4NSVxfyBKWG9+WuA1iXjHQrKlLA5OlzR+aZXQkI
7F4RtrhSlwO84Zmpy/ddOfoo2E6Zuf+o8XFibxUPWMY3GMuLGZvVeBoC5puOfZj2lQWScPC+p+TO
eQ7SxxCD3nAILg1TscwVIXdcvIM/5jRZHtnHkwWUVdxbd/NWcOOBfvMmN/mWDHCGNxS4t6NPgE33
bvGpIsEIcI8Mc1oyXvyzrKN+Xp8eWoLcp7qAl+JT9p2M9+vp8wU5b1WtGDlNtDQTAbkalT7GX356
x4jxfqHo/lI6pfUDp3qArum4soscmgEOiR+illOA2R0rEI3Dp1UkcphTm5JAPpFkNI5nBnyvnSK+
B0b9Uicmvq7V0IDxXvcpFfxIGiqYMwD29GCAx2WGCkOw32EEkwe8cXNXuPfQk23SiaIJzQHzGpRl
yPFcUfVEPZCUUxm0jwC89KeI21RuOrMTO3dazHMAXXSzTNTnf/VQ2LtvfxzBdoRVgD/axaTFMa2s
3rMnw2jrAIRZiRaIo5XpFf3wzCwS33Bhh3x7Z6ssD90AiUPc/sAp3CdQM/O4/SkWf8W3liG+BFEP
QZSAXCNjw0B1j8Me4iVxJi1GKA9sE9Ih6Ekm6N41hcvvsBh+gqZvIZc80+7+QCq6tGyeIQXrgDg4
ZEGffd+937gpgRe71sm3p/CuPfhqk9adOLrMKV2KvTA4XKZtUJk0r5EGn4/ELeVNPtckePIrm21p
qmrzyxHJzsBUoTjU1llKAmBndb7GshSTpseiuXUbw1wC1CpiFwtghe5nY+1p7mrXAYIN8xP/ff10
ueXFd7/zjH1142Bmprl9PnRGfrbaA3p1AN5faD6+dNBoNcCj54lU6XyUEftTw3uLjB4k7NwoPJik
tszhj1VGp5o50Cw85r15YWAbOTOGyvxEN460AVwQsJvTklAxxAfpu5SfkmKr+oSEqsYevcKUVtxD
5I716rtR4C944PxNA+taaibrHxeosg3HLjAsM7wZo7QodObb7YSdbQ3lPZRNtmupwlzKlYDQTnkC
onHcyU3BkcFuMk50biNPVJiZR0zv+3lV1TXO1/ILa2luCdaAlYD6DMxcJ/UZ1bfnVM2D/Tp0c5CC
xXwxTUn55KNRQn1GEOCElUfTIEIAHT1LBbOOiUm+x2QqsaSZH3nsVZ/fytN+TWd+LZtQKfj6sYQN
M9VRP9+lITkWZ4h3l2Fmn7HET79dBfbsxOs/xU5qyyDtvuXMv3SUSph4k3GlGpp08W4NY3pFsiT9
ikWqHl6hlhn8/r9QuXLDesR4KZXx6l5xBU6BMFr1FLvSzrmaSnV+NVSTfQLaA39zgCFeoiIi9IEb
LNQpijRVzMvOimjsbAF0f7uoCNaodycfV7YuA2u0lA4OV1+mADBQm1ZaX62XM8tF7qAWxK0mNBiP
poYVJee1kBbpLbIBqMFVCVSXnU0mu7AK9mozMWkokBCgqUW2ZB9++6Rz0sLe84v+S7uB+t/6/sny
s8K+oE8kD3nhwTOa3g/yIu53yDDHDND2REgaCwsuMykc9178lLPUduXBNImfa4kgyDfHAMXsnGhB
mKPohRynhUgvQUGyjVlV1exNxcEBT1fMf1Yc/0yZsNRR0iEvOHcHPBu29yhmTLYzTnGPYnFq6ojF
N2evfIZoeeQq1GJwvvhlz0YK5UFvLq34mFOoyNdTlpczhFbfFEkG6j6c+1Of0Sj9NRT9RPosU0Qz
35h6Immy4bQmKOPH4dAycMAkcOk2ECMpzuxGM5XPA7lFwCUJeDJYzAzdB5UTZ/dJXBPG9XoT5+Xc
438/jEmVtWOuF3j6sZCH9jTD1yVnE+IPaqP8Y+0L9TZ7CMn4G8siGTkp+BWJZOfLmETIEVgzDBFQ
l6zDDymD9/Jph14xNGTlGqr6qsQFq0EWMJEIbWzcVo4DekC4gi7HT8KVmqe5YnI2nsvJinpli8GW
ZiIqsELK/u/j2qSGCepUHt6E+ncwlgRwNzrSzdBO7B+GvAGyaFcZZuKRc8U1iSWWWCqU+VcgMeQa
n3p3DAplsgk2nemLtDfSnx9fngEsjZh5cAZ4wXKnaxtp9GI2YRZjWs4lDnNFM7zZq577k8WIvP7A
L1Ej7Gehw4a7ZEi9cilAOtLNeHIpcUCv4ZI4VfrVeZ3ig6sk99maylmsXUHbaVmxSJT2TYJ+Pm/F
wGv2ijB/LKpdHlrvMOU1MGdJQ42b/vYvF4aj2fgvAQsZ18aLTrDs0MRu5S2EBQWz6HDe+OrABr+9
CuqCDL/x42tP23HRiRnejec+Z6XeJihiLQQsRUJjd7XAKbf1euwN16b/nZ2skgPlj9Y14OtraVeW
9yYVo2mN7ijJuoHjtn7RXoUCZHPogypPGFirw+82ldXJoAYLir1BLTYV8uBLWJ+oJBj0HIrhfKXA
NovCMunwMwy8rdNz+EuPDuoUNF4I2j4fplXwRhNdVOKQdXUseturDcg8b/Z/E1M2PEsQTkI1Zj+C
lu5MvfHcmTwsoXTO7Iq1iDISBFAGamaWJ0ixoYlqmhcC+m4q/FgVlao4E3BLEOGj/BCUOazNlubr
sjvACi0uDtHSq58ju4KLK1rlfNNkfqmCJoxhcS2KQ1FUOJV2KwI/6hlZfRyOvaq70xgR+fQF0tZ0
TvQvQuO9M5kcAPiL4RZJ4eIVyKsPmX6qplzE/oclWPobgPiwfeOpF7ylVi6ufv4Y7+FC+LfBfPED
HLtCBP8TR/5eUmXZ8BiEj1xWxKeI7UaAD789Xi1+HYm2IWgP0lhL23IOrRUVqMUuqfQbVBYQKim8
O6F/7MKNhC/4Ybq83yMhnFqMROmB8ySw4xwzBHxM1DT1NAJ9EZIuyQr1JIKn89stHpO4Ij3sNqay
+7vjGRVZ+WYzs0bEcijtFYjy7rv5TRuOij8Gn4XJGCj4Ih7PZMLeGfXoxAY8Mg2ve+Qzm9T09O0o
9HTUnORwYgrwgoEdUkCGZP6FlHJzA27HnNEaVTmC4RifxntxL1YcJ6KY7EHm23yreRFODFCqTFOh
51yNkKCVyUc0GSeaPAsZljV9iL47ZPsYaMdU6YIBgyony4U6io/N0rFImP4/S2vGwrxnKQbLTs01
NDUOjB/GIPDh99klfML3zJEmXwmmmWJq5Z/RaxN0fC/G6W34f98JBtb073gpPjdGa6wrx+Kw5l22
7tia6x8b++Cjkhlyf+gkPDmMU022jFMVF9o4XYSlNwO54WCLxNkLKNRFR6OjdLqjhHnoiwqDSjhp
GHVVnOyI07RuJbxP/e00wp10AT18jzGPrczpcncK9SS5zLhHk/HQa56JLsoVUMAfBHpsKLTHFInW
cLpvunSHjzkp+TmjMoRwVAZx6iL3W0JaqyRMdFpkT7YknWKMFuIfsZZbzGKwraFahowuOmQfM8If
siWyXSAHzjF0LAY7KkUMYtx2uWH0OkLJ5jn+4XYijKQt1QzAysyvERH5CzWaBF61dOtdZV1b5R1I
3hUNu6bISA5hEluP30BayaInlB2ZzRwy6lBguXTFNdYRKjqHQ/47KiGW8SQUPVd6TWXmQS8CiHbB
+FPDLkxVefB8702t28e8pXQ4MogZFS8ngV/Lj5Vv0t4pkTN3Inw8/IHWRlQYrx8KYW2f9BVtgMBU
EarNkDwyWtkd6Owm5KG86kQ3py6bta8EixEcK3Q3i7WtpI+jiT/dHj/ilRxAL5IlaTtjWWLt5Phd
gsBtHWqO3TKtXQalmu8afdBD9VhIZwcEQwP576u/P3GxsJGQXvHmMUwegu/LOn8VzDrssTuAh0rC
7FiUlIMYfal9RHp+1vuzMX+N016xz6tkQXMP/vDArXoBRK7gNkba025y7b7V+IhUX/4PBm9IZvR3
GBhr6wmwQcnr5c50nA6PATGnsPNYZ+DPhSK5R/z72I1jyShBM8zTyopAUanF59JiwW+dvrGbrZjU
y46SlDYmXW7EAmvJrQGefQnKx1qBz+2IEVOCrIxOeXdDwB+ei5G4Y15f/OFrYAVju9xX1oNzjjVW
hqZZkhZWwtDx1HkSOEXtEs0hZ1lav0IkBcsBZtrB+A3zKJ0kQEHH3WE+lO97uqgONcE2J/3UYVwf
qSp1XHX3vW9/ftBWeH3+pk1CvszwuWNQOT3BDqVJGRAYzzAt+bg0oXQb0NmgHIr4rnEOhHQaVY4A
386HAEbH+6lUFMB3QKySNyWJPRD1Tvbc/EllO3zpDzyDuD9KvtOnM4Z6AVXXrqG7CiPEnBoTE8Es
mYTaaDTYhCHWGluXgrSlahNnUjkeqp4bCN8RTkS+VdcHluADWuSL21l3YzF8FRYzZyze4HJeyxdU
esddQ8444k+vBofmEUJfRiek6b2LAh9aldys1VlDepRn10I6bC6gcxlbl4aGCHhRUN0ONBQ6sob5
cGCfbTmZaAwi9qoljFabrMWNz7013xfWs3/z5qlbLLCTq9YFI8Una3TJ86F/1jxJj48WsdMDN5ab
g4m9uwVxEJT4xlUc7vN6ettiSrlLHIhZIYCMjNYlMfbVvTrOQXIpaiCtF7JPxTwDSDQ7D8yMvo1g
BcnGhV2woVRI378XkNeYqILVWSngysprQwqCbjKBiS6Cj3vWu4XhJNeQr1LVN3b8MkrKx2G3W70T
m1UYKLf8n9j9+MfYAFVmHUzKTC6xi2e9S3bZOC+SWWF88sdM2cr1WhK1MUSIDaoXzEUaxXUk5zyu
Kh2vX4302S3OlS4vkFcv3Km1JhNGnLYFCbybg5PKBxa8wsYkcNTH1WoHZqEUbuS4RbIkXkQb6Q9b
1rLvdIq4QXbPTmymNWXtO7kwIm/GlKndsWJq1xPeuTDBh30UCPv9oLLi1Q0pvoMsvqjN7lKXFZ97
goJiZxc+h8G7ujs07kbHCSg7ZaGzqo83gyoiM8tka5BH8lrUT14IPWv7Dv+bVZoXud8ej2vtqpSL
fqblbp24fQ22w/h0Sz0gj/ZMn8hHL4x43oI6kuEBobTIK8oHPir1yOOcPjPAMtz5Qv6CWQ9UAuGC
JCxnZ0QX5FjAf85T1wA4+3rpQNRCAnhmWrk8n2zlDyVG9Z21fuC+6A2PlaKLqNTvUf5D/bGf+ruj
2QOziuEF5FLh3mAVerG1gBMW2KjNCQHh+sVsVWSRvS0cMFt8p4HWQbRbVpJ2Q8jHDcMm7jkf0a3E
pvBSMACYH7MoNth8NDC97m8c2BYFNuhUJI7GODVFdvdNGRgMosZWDBY1Mxd5Ql4NWZ/Td69VuVI6
6U/MA+LrOubnhBEzEk0jkupYmFoXmRmG0HvG7MuErlrc4cdlaGguTQWdWLK+re4+g1qxiiHFRQMm
8Rf0BpueQ8QyPDe+DJwIuDb3zyApoxNtSLus1knxLtFr5Ang8Z2CMGE3sBrueFfVNEFovQkNH0HU
7oI46buOf4J8HbndEqzOd57DpIYreLLAyv6Ket7Ups3bwQKk9tcIw9F93i56wBl+K/kl7pfYNH61
lW31iQ+qRs9rGqQKXlyVAvyRiQioIb38LgF0U9pjawZl9zDnpuyT3zlcHNkStuozAJ0r6wIXHm3B
o3LrrdEk5WQ/mV4qREdW5lTHDYSHHSBk0ISyayX7JXv7qxFNgWiQHcFfdjYlO5FOmezQ9lXeSTpW
yjL/wTZtFhMhDnj2zgJJhzKiumNXlaG0h4HeymHsa024lze9MdsmmJLLocHBYeP5nAVajt2rU82s
VBYce5q5qPn/3S9L+kwnvoK8/mB9haTeQbbTCj5jemti7cS2gsPG/FLHS0a1/fvcsABsMd7MkuWm
15pkeAk5ddk/A+NQj558wMGt/dfuDsWUiufWvTy6LlUaEfZlTxUtrCW5Qx0/utCOwUQy5RkkRRhL
YkB+61Ox8KO9FG2pDPYo+gbhl1SXtcQIqqQsDujP43goObrJ+kkmBrAwtZf39p8DvcfnmAu4pWYL
5NAP8iFFnA7OSp0Iynj6Zeq8P9LBoM2bceEcarzHdiZ1Iw4H4VKS7TEDHkp1eOViPahq4cJoCFtz
Fw9IPEVsKIZ3MH8zvuMm0OBC8BDhUeAtQSIuCQV0hp+NLp/wb4so8Y/wEV4At30y/7a8iVfsYWue
OaoevzpHpLqG2xdEnDNZHUUweSRDcItER6sX1e3lWSDceF0BQcptGpQD4M4047Rws5oXuAXLE5Mh
zYB2ZvbLMFgakzO3PPav8wWisirGSOla/366dm5uotyIs6GV5g/P1a3K3x+NF2wYQl7Ue+6uBJ7m
XkEdDyVKagIQhlFtYNx1eY8JlN3dTFojtWMu3lrT10x5fOFVixrdRxFV4r6u3K5J7CyPlLOdGJuE
5/ZHsayKuQqvqcxrCbzK5UlBDxu2AIVQjf4t/en0X1dwpSR1vWV+raeD9hehdFrGIjPTjWyAqzGp
0EjfRIo6ovUmPzQqQuFFacEFk48o8AUqGMcSQNrqhHnSfNCLSjNrVtbofT9MzvxtlFAIL6LrEN4t
4TjLhc+KczjJy9sQY1anwiQiKe/h+3s6jeaGqp9EWiP0PObipkPaS9689ElJb+LJyeZTgJecowIg
wMOEsedZKyn3U92zUatrltZPbELEmzRU0NpWGFMKiwGp0n9xdKy/Q8qbof7sOAISjCa6ys0HcM0y
f6+fypdKFIFIpKxSqeudKMeGtAFEE5KbQNeQ0xwFrknyeTp8aFpS8/OiRGR28d3yxNblbWzJfqM0
Y9FHUQMfYddlKn9CNgJUyq+FnLMG+QOXDWhvwTirKm/TXfbTVn65ZT/MpnGt+nLPnITB8GY1d6wR
kBwkKFBdPTMasLKGzLiTc76dD/K5aa592K17GUmWu6VYrh4ZAqGA4U3TwVW4jxwzbwtvJXJR3iYh
l4FJwjQUxMS6MrzpxROaer25nNX3jjYireZawMq1DIOe0IzDM9JLQVK6ELr+/JDzpe99AGSb8eFR
Is4TGsBElg28Nz/WxqhuJRFRvtV0FBQPM1YsWkfkKrycrSCJjVU93hTxu2HYe5pflkTQhIPoVNqn
T3bOyqf0nsrjd4peUZlFnfPine3ycZU8I3EvKAo+BfOAI/P2ElNxhmWk8r+9uejTRhPQ+guitLWh
ZJhRvampg+Zb4oLQDUQLrTOaxG3WcmQmhsF9rfh8wZPclFeEF8PZfC06Jmy1CeLJbcadNnx3fBB1
4vVAxMNSgUcC+ZcelkO0DNSCX2kyHmM2aHRsJZWsnkmoHLhevtqADRiOvIwfXX3e6judVF8Dvk4G
4hJVyCQEh7dkRrISSZKevBtxEG2bPUEYQUupnXAobPTN5t8by1NQtf0UlhYbkV/zIwu/5TdK00N2
loqbhaah4hckompiP7s0XpLGbFhdVW1/s1I53ZkkMSdEzQ+Nu/7RJDgF022RBwlBGP3/QKoVM32p
Ch6mqWdnQrekJQ3bFD3mqWFhkLSgnJfPKuRZU16EdYIKxCMj2bH9QEcnmspd537lRyzI1vPNjzWw
2mcdBtf3M67huCp6mg9ecjfjYMxKkNRZaQ1riQ3hl6iD5c/TSPITWlpItKmuqlIQ9RPpgAmYCNMG
7atf9S6X/MHzOrnHwkbd3V1RFr+NxvLSR1SIxiNi4AeZwKlOUAGelrEYavJ/YpdqjDDmHB59MHNP
lLX5+MjO0YIyHnhqmhRw98xfeF1ydUgjwFCj3gATQfQZYiW6wsa0ChsPq86kmuXz0YlBpDpRPNz1
MHOTbEsoiLW06FmNvdB+1STWizBIbvvT9fE7wZQFA/ncutSnZhDctDeqzcfhMX7vEZQN/k03nW9e
R/Thm/8ltZgrl7VfJDMrkLy31S2Ui99qbPSU4vMBcb36mBoXjfPND46hgkj5CBmRNTBP0ekCq4fV
1nJrO9ImW3nnBw68VGv5IEWcXkt2ujT0ZVfG7/bGnINiBaCDW7e15Ch4nsYcuB8VIYfRGEFRFN2d
QFGXlT6bvcgSB1W0CfISpyUlqbXxAQUZyiTX/fDdkeYDpfKVqQnZ27z9bSGr3umdgDzCfxmQb2Ql
6MgkEkxfAo6awleB8fXj65XgkRvV8USCN6hI8zs1qy6gX78kmHO/+4G1vQntNpJgY2nA5DRIXxYi
+i0VfwopLwINlsppsu8dNyBkITB1/MO7WL9uwC8Y2dnxnuwNU0ug2OYp0S2fExzf3L/QTWf3D3mG
xEzOUl4Ey4gqngWB5JXyeKYnV50Z7m+8lf9DA4hQNxr5qFWehXu0PObCa9bMQcR2zy2+woP5MpX5
T3rghzkHjlRVqGrfE+P3a7xTfYRRtGMn37cYQ8Ips9ebX7aZBDn+KA8wdr/NrikbGLE9hZEulbVS
T75emfM8FpTPrxBy/U02Oz+ko7c6T1SYPBUTHlh9jPa6cciEj59sSdfbRqTPawP/9kLHKA6LESj7
ZCVqCNYgTLRDJyo3/w9zwGme5ZeuKFPxPnB4GYy2NHnnBFrnzN0m8uQUxn3XJrTtLfhFs/sVhiyp
r6I2yYNemTYOwkA7+L+dJvOnhVdEyZYW9CL8+7MfXh5HXTnul/ydTls/M5tgAXF6K0CC8peFKSME
CQeFvDLqdFM07q6H9TSc9Xu7Ycow5ZUd3gzFAe5uwqYCOZmmi7cU6DkS0mKO4tmc9zf1cgcVTFaT
+mq0TxU3Gudim9IB58c+yCOtFXeoIgKka7NUNRFZBItK/WEUPy2xvHrXUrpET3Yl8T+xCsyrE/Cc
SyMTSK2I4ARHKGScbs3VbPyBVfpy6r6XI5e5XfcYsOYXOAWnFsq4dB9IIKzXRIzXk/MIKvJnhkh7
HOK5ZT77J0O5JiFIPc3JHaX7Ojqeri+m0RbfE0Hgnp5mcsVwnw8zcqVhXhqEcz2Eg9nDL2jimjPd
fu9C2gK/3p9xpZ41pzOSNbJbBUfld+iRT+9kJOjdx5gcuVWYclfyW9SamCg2AdWVV/bE/Kl4DH36
Cy9517i8eZzqySQYWD2hFM3Znv17Vw2bTmU1aOTskrg3Vjb1Ml83GSEC21QynujLxzfyrvjAWC+B
qelE2L4fLAsGH6MPZx+PX/wyChBkpDsrejz8Vjc2cNCP3mEGKadh9nwPzxtxYaAis/gTqi3nzKMT
CXPxTHpt6kMjqC+JYa7sDIJgejcnQ4LDQe1y4dNXKGA4wWIGSEJuAFT7VfBTTLSBf2yI7dozNnzT
u001jXfgcdymcYEqJ625Rv49UyvrqGI1pjreIIcmx7D+6Csh+aoxkFuujylZJjNKbljT1z04e6O0
nQDS/iQ1SZ+OayzSDTz9/ZP2ADEYFl0Tfg/TBbrUgJOJbRxhwTw7omps//Dy9yo1UYr99od1ULlZ
IBMPnhZPsA7OFMEFXupZS1cAP+rEJZwv+tFkm6ETjQh9aUZe1QpoX+MMMHH0usc8v+URNyaAfViJ
cU9m3wqwECXChOJCwgWVHc6TQE1sgN3QQcHf10BDh6d3KtqE6pf1CPHFbzu8dn7L7i6qx8znXzOA
uwpU34Lh9g760B6j5YB1UAwawxtAIHbsvalANBFamrLOSzv2WDkUaTRbaNhMZjcQ1R82TYjgeU9z
6fRbaWAlbOE/l6h7rK+urCnCTJDCr4mZWUL0QwhKjpdSjM85k3x7At+rDjtu/k1xy7dL2Hlc9cKo
G1xYlgk3s0gyl92slq4xBU3ZG+ShFZ0DVljjj77EAfHsPWArU2/7KvEtjF9vdqBuPC/P1EjMsRs/
SzJwdBSz0hy/AfghUiOE6xB4ucZkT/4bEHNERcq3Fcdi6QHeZdE7o9iM3q9b0bM9QTLFXjiWhg4H
II6V6l02OY6ng7YmW9cvou4p3qwkA2BEGVJK6DgPE+gX+flpFuijApMtr6L+8NejEEJgzXRPJ44t
JUHZ71DhaW7R9SpBwY663SlR+j3ycrxxmp99WKtbNANkT/tZ+LaZaAZbttJnhLW23PkVHPMGY422
nj3KEyxkv1AeyBRjPdXZy62A1DUEYtwQcGQzwCR8YHAlH0nER3Dr1zovJWDv0wDs1fZq9S4sUgEK
W+qjsWUeAeIyUV2navUrGocKRbfOUfo5MCR+fzWNPu3J85ToMA3KFAzABzmbbs4vaorF0/XDdzPv
GI9UHEoEXIsypEfmGQYakeKG+IeDS1CZ+uGe0UyZeMjDf5goAyQOl5hUHhnl+h9qfcThgXJNIX4P
L/B9dKnA5kYs4cfbSUHLU/sZ12tzr8lmpWq484marQhphjMRsce6EvFUm2tX5EZxwtEZy/OLUAp/
5pBQO4cfwsuY3s994YrjQgVyKZSt7B+27Ci7RqBDCgHATwSC8ejgSFnJRHB5l3avpAFida2biEVR
jsOfDfQh8CrgrfeiZ5/oVNShbLfCL1wZPxPY2DCG21rip9ZWq+UVSQoDZTEqfBLTmx4gGbkURy6l
pe4KfwhYkVmEp5kwCQx07mHetfi5z/9vpUP6tvpQvS5+Z4N+b8F1Elm4cO4ofetINu7ETJKf+c5L
HUzTJDtTjPomYI4j04l+GIwyq9nO23VytaIru9nwe+mLGzgBLRMFJQ5CUfnN/aCdzuLC4VoY6I6I
OOR1slX1m5Y4ujiCENQwun4yf7LByMyw+YcKv+PXH4XqQvN/2b02dU+mcI1wfPhdStmhtyXBNEN3
2PZ/S+RBmHjGTov4sRpus4bKoWz6F87yoLFzijAt20eF9MKpAydKI3YBaAAqWPTNaTk+Hc1Jv4JC
WK5H1uEhfUPC6gwbUi7jjCcPRa0WK1biQqg4snqroVvXYixD9SbWhDrSxvhGvXZQy0+ONTbNe+Lw
Q2teyh0ux9tt2afK6+51LlASMs3AU7LR3VvQl753FTWENCSrQviIAP8i7lnFnOIM83Za+JAJ10Ii
R2Gg0yDVyhYFG6jYqMx+AjZ3dtinf4tpJ2rAFA8NgIbhkT3ZwtouEEawHCwkJ5bx/XqI4eH6mVwt
X/jLTtT8cri/MFibYe+Wabo1iJ09JCOLfn6RpFKbKPDS9FcWeCGaSaa4Yc5NZtEFJltDXxLRkS7F
JAwxhBT56+XShF/DLPR3ryQ3lGsMp1aImexqU0aipNr16mknLGE2IARAIK6e4JnD/KVmRozb/W7V
UI730vDlLjkyc2tuwLoYV2RFXgFlFa3uYbTkFp7XoBrD19wVV9IuwrEurOgyqlUqOb226tJ3rmiV
ChucEGUhUlZXxYMFWwbfIotZl8zsCI2AD6IfL7kRcDjQxHmCPGfRI+haAJEfjuYBgBzVPW/U/lAi
T7Ws29X3h3ift0Ou/XhkdXOlE8oYs+/3I//Vdp2haA6GKwdvfSo00zjpFUU6kuo4i0KqBw2wfLm4
L7GymQlt2AuHhiWhRLLpwj7cr5t1G7qQgMoaqozNZ/lEPX0FkTuoX2wihc4VtWNzevnPyZSGuOop
joJoLwZADYI3H6os0uThclELUfSoNBksmJaQCmNIk4KYfN/g9yfFY+Q205QZ0CP+46MOufs2NQNF
iEI6DWDfu/AFq8y6hNgCNL2RXmv3mRMPc8R01/6CVdK5/FPzzIW9DXXkNhodvw8TGtCSt9iV/TSW
TNVZqAHmEezz7pOzjNBrtYAuTv4ykYeZytOQLUHPoM7085JL1uj4aEQ563FbjHTUQNqv9bUztMY/
6nBapbHQpAmSobLuySGEdCJ2vqGgwvlAbJRRkgEwHCUZdx4/nx7YnI2DQH7rdtKhO7iDlh6ta1Yp
78DEgDccWV0nHz+gM/NzAqvnbcD6NuPtnYoSLoVFGZ0IzMR7ESOCeRklDi8/hheutR4DAYB1qz+o
lMnV9+zvvgwQwTx7fqDo7Ujl1BmQrOPdtd7Z49PSY7XRuveUiUfD7NlwX3NU+SSi0Be/tvFpB6lO
UO0KPH6JGI/T194ipn/xsukTT16k6lM1pL+VdaONRwRSQUFD8JIg8TkpryY3dLZ/66jhJXVSm2mS
zLsIICoq5EqdEtkSW+sm/4nq/ykg+dykli/CuCp9Jaxivmt5TYPI5EjLFAUoi90mmQSuMB1is1A7
0RCmSzSheyzzHHIuBw1WFIlm8pcMhXzubthItdX/J9jywOp45CwNdTexMhPq3CYOEOikEHpH3M7O
qxR6jnSscy1J2bjdGz/p4FPi1pyINCzCDX5IttrDX7H1gRWMS2838N6LNLi/uezszh+vP1m6bX8p
su8fNjHMeYJHnOWp/2QGo08JLnPo2dlZ5tyyrxBWE9C9DNgKK6+yPuX6YYBOxHz0GkfCp0nYdlhU
zjr8hT8bVGZk1djjvB1Yn51sjvTuY8ZhmfnaKla9dqwHE39muTSAWcAvFdPxd5iEnsfV3+6E/9iH
W0ia3Us0qCkD/GgHJWek0zvFHAcLVG+eGhdq1wg+MfIBqlKGDgBHsMPR0xwEbOurjp8c6klPWCMp
YixP2hP6O5dvphfcQytV4l/SYoYA7MY+QL02WXEUD8/QCLBn+9F1FHCCht8ojiaZKL5X3OSDCIcG
JFmf0NQKlWNlbaGqC68c5GVLmCo2OOVDyEDM62TbnfMeHFwjTi9w4lcfEJUIqfCIVOVwDqbBs5G1
AWbNzced/g7VwmHGOtxyZVMfxlennroihxOrOrzqUFQW1V0JQwvBWgYmKhCdENYqvCOc2I17fa4d
2J8sayncdqmVJJ/OD7eLOLkhaZg8ZhM6AAzPUtWAMYZOAHsNwpVVIhynRBSX2/lgWQ8fEbG02haV
NUWXQYOOGGEunlFzKragrLhSZRBhDXvRXqKZU4FDmUZDTxYNkfqYeH+VFUkF9mCJdb3M7rbFNf+5
xMHbFgDQkb3KlKD8ign1esLk0O5eJzVuY/w31XDnUEbdn1f5ACLyUNGh//RaGAnw4l6aTWcV4tIT
7z7Wmz/F7JsG2kE+6mpcI+ruyFo89GCdciYc7J2cHWZeQ2Ff/cyZ6ajNTqP3WvWvhrPcpsGDNa2Z
IXjKQgDA8g5oRbxzpqxnQeysS7PAsit3JojBd5cF6wJkHk8bl7mbiaT24xpZQSWQbvzd2i298T5q
rNDm2jD33eQyMwtikSGcbGXK+aYQZagxyxsc3kCYKdgulcIvVfX60U/Bm0AmvD5cGuaPd9JVoe4e
C2zc5JKHSeIfR2xWXGlIqVafrbmacMbac4xR/3uEWCMvex0YPJRkExZ5r0ztbG7Mu+Pj3GwuX23l
0U/fc1ggy6qD7qUTNgH8G3phOSCsKx7ufJC5Exs1CPDcU0EHVwkTnlywGidTnZbM6K2hRJ0QY1a/
ieuWWxFIz3k9lWnF5EySXeAlY0AzFFRjASjwupGz7GVrL/Z6PV5TeG5s5qCAN2e5oyjMKGP6E1AN
Bw+Ju9gX9ugL/2jfnuDNAUpCBmbZKi501OtrJsXuoRhwbqm8cBTxW5dLPm9aNPrQWkoCq2p+PG3r
fcSunZTFCiN1CnxXe2KF4hAzOTt8PM7iW+rM56oi2MrKA4KaHoZP1WiooDR7nHRKmI7OKh/nkGCC
nUiXDKQkpDUFGQSyCsA2jB/sjWeSIBhqPxDliReA7nutZaFNr/e75Y1tKefMwof86iNR+AzaORsF
JWniwocLeZNKDO4jKJSXIZlZKN9G5LI+cV2Sf7m7DhdS8AAXXNkZFSdo2S9n3Qv0j74eRG3BT/fa
Vdcr40iUb1FlDfMmvHaPW+6rPcbmSjQfCMMysyHCiSbISAqX2V/guKK7ZBPRs7JOvn/uDJ9N/5YK
ETh7QsfgLOXf7R9qBesby4NeHyvOrK4ZaVPA5U9yin+VlCrLALLpFl/oPGmb8P6QgHcopTe09JBX
68T4nyp3NeHqwcLj1k7a2GedT/inTybfaYvxxhg79May6TDgsZjaiBBegt48GJZZRcqiANUbF4fr
feP7J4TSZ6aC5Ufvyf0DW/Qyk0j8nZmQWu5rkrUBtdi+qO/NAjLQ+6PtrCWLI8iY6vlfdwflVQbk
o8iCkQpqCljQG2xOpWF7l50aJwaWTBcyerUqXs7P35Bgcc3i+QXshI3N3/PXtTI5Moy8TN4uXqBM
145R/p/a27/Ql4PCRdKY58sSIOg2R4EXsu+AF3cBOO5mYBKfwwmCbFVMaYdJcP+zy6ye2YN6M6K/
JlEqLEXg5Hi+dcovc2QrBKeeNaz3YxwEh2XX13PrePs7UuBdD830xFdLxBkWXPes9n7Ty3ibAABV
oNNmhYfyUxG8zWJJYrOQ+ExWHTIJBazxfpRZI3DGjZmBsTPgHH6sACLB7KrmRgDjNoM866Et0NGL
lrh3NMoGRu3lg7mA4j7SZEr9OQJ8X6+MkwRp0RYr8+zrysU9LPEXhBYxHUeo1mO0JolDyotneg0v
GYhqU6luO5WelJf36zYe2iu3eOTTZ6G0M4YJDplKwiaNafReIUJByU9VmIfRcueAxo/gcdpC+ps+
Nd+xPcfopOqwggiJAzyvl5qSqNBt4XdBMPjBUJ/8I4wnYYwAEFswA7g8GumrBbxMyEliT0r+lwkp
dqqg1VYqCp2o6oBtDiXPYxT7IT9KtthMwuBpY50S41yPB7nEUwE3OM4BXrW/xUQOg7MjrwxhYBLf
VWPImQyV9LTiKclkLBFzFtFo9+UP+DT7nqjQKZMpAfen8NW1hH1tTC47/rn313GPBgKjgwU3Bx1z
whWKl8SL59Ucp6QazgAuXxc2nZwGLkoXiPtLysP1VlwRWkWwUmGlmn/A8QgrU3dcP/VSDIJsYjIm
sKrKqd/q6Y1er9EcIzL4FR2RLaf6tuv9VKVwpJ4I+4Yh0ilSmvTnG1w4iMzgLAOfwKmotPj9KtK0
t7zKJ1YE2hwsHUKRgzLD1Mwxm1zMvpIIZahtA7H5YJw+gf6RkMGQ1FDRYX2/AWRAD3rBaozDS+4X
AzCTHVsqkXwNsbiwEV3Wyzv/bVbTH6UzgoTIoRo6Fy0m2Xysd0Vz2mYKYYgtxjsiKDiu2ExQGjPK
3a4GuW3rEv6mdW4kK6TuKX/kLGN6lVmOeQmRFY41y8IfnjudJ/VJ8dsWQc8NeawsU9yrmEYzYbru
xFLk2y8rNlnMXW+sj1+e2pAIS6FdzJOYSfVflyxC5d+oYVW+TOCXm3pwNU8mTs+I43CVg6a+vRg2
jEaTxwBXA8QSMfnTYfpSFFQ8aB+QTn02H0Q+pfkJ6Xy0o4Pq8yyVHA7T/3LvRC2BAqSe02HTpjNW
/S0w0IMHBds6onRXHfcpyOuQ37FOVp7KLys7jihRNWFSQTnjhcOtm5MTZw+01ErhsjhhA3SalTwP
QlDd3OSK/ZC5DXTRejsP7tDQ7dmWvVeCWt8YashAfWhaY17JCIJiUQdzdrf+dIpt/BAndd/O1gEn
FlF5B2X40a7ukwhHAr8Vw1l9JLBomMIOs5HqB4lPud5JiIx3jpVbfC8p/3Q9rqamPt+Bnq3AZiyp
vOFcFgZ/V2L3fZnPSCO1NNj7FuQ+h9lVWn2EgPlWu4dY/fdTCayPlL5QaNeAtSNVN7yybdEuDyw6
7MBBD1tx3d2OLcTzUOX9fEyoaGfQPrJTEcJtkGS/2/SdqLJPjRFiOgAP70aV8zrBkv/D9AF3/fVJ
sTddXhxb7Kl9WX2U+7sClMSqYStkY86qVj/J/fuGvoCix8lM+sPjGczEGZ4e44Aed4yIWEaTY0H/
nMT+yUO8vQlCe1rWwUZIuqdJ7qnrJ5pa06tFQZyd54Rd0orPDCcbfRptpzLUHMwpIlju4DP7XcbX
zPU+fTdfoVbJGXL6xFpqKFrunUCrLFLxbg4fok+ty338woRwGxXE8z/WZ/OdLk09IW+lMaiMOka9
vzu1c2ATo7o58da3UFwpGSyiIT7Vgql9My9sDINDhLtOPIKN3A5i+IP+eJV5rctjctFDyuBeSt6f
EeQk3en6ctc7cZe9h9z/4ZfpEm70tAuLm/8c6t/q6XEF2XoMQUNCaO4DT5i/4xv37CUsHYNuEk/z
55E3rtg3NwN67oFrch/5/D6fnH9LB1dxVv7e7Uimmk+C6QXb0NeQOC9q/lN1uHsu1vsAr4Ixd7HW
VcD/hy4nnRaoEax8tjUzcXR5lBMa6Tonl/svSAx0giYLWAIxViDBQ76/NpOWKbZrGUw2rkVRCuhB
zzKhAjA0wJ2luKNq4ngVXOHf7BxoE4sio2Q0YGwr9WBsee0On5U0G4F5azXp2fV0RGEQuFjxDF+o
pWr8o1I6O39gOaaZ7tzsh/p/XEQLCADFiVX2bkDQnYJQQV96ysgjLksrjL31NPgt9vebSbpTfO7I
/g+DkYiG2Ul1Ob72IDo+aUE62nHHEFhKdMKGW2b9JRGewHwpAWdslEIOmTEANJojpvp0evPOkQ8i
XlhBkdCtLIuqZlxAd+CBIuG+ivs7qcPQnzUZ3yE9q0f5aYNPVMAvvzzXEqD47MP74cgooQQrKiyC
YdMCvX99Mv5k9SUzq1pXXZrlfjJx+TnLDa53dVEw3cveSd13RXjTlkX8pSB+FYXKUCQnaqzb/jW8
9hiZeRXvChokl9X71rhtjkay54sP/XJMbbsABun3kAL4OwiQUS7pXTe83K9odxcw+qhSv6UX2svH
abNCta0neGRV6dp+ah2M4JZQIMOamGF9yLGtjInbPy9WbDWUpdQk6/HKZJbpyzE5+0/heWb3hzTk
vRWMW+w802eRwAE8yld2l/Clc5avQ0DJOAg7whBwCtyJykvROPqj86kJWcaY+AAHTONuLxaFbipe
KP5dewUaAH/8GiprTcsRcHzHaTuEqEc8qiphx8zsdrKoIbmAH/rPk6H7g7QtRwLa6amoLwmsHnum
CFKEPALz2WJLcIUNs4D7cjH7cjDUCxCEi+ktSXc/mPW0Oc2CmuqkJZor0RpN/ZUtVk01Rgf4lBpg
yVwQjKEhcbueNitn6fa+WDQPYmGN5kKozKotU8FysV5RuWqsxNHmRpXwKnIqYuzpLMhfAevnL8XF
P5cQZWPhAoutkkCi2iQqdYuz18Zo+6UKav+ew5pcEfJwjs37LkttTwP0Z6oucsXgwejB0cffV07k
0w4f0i1KAb4Krdy4zxa8ehn3+Hz/b6rr2ip/hpG6MPLggh8Xg/+bzQKPi2IlyDpjhN+txUwWY84j
ii55HwmsqcnxbdlCiHbEQjZ0etl/bPX1deNWQbmc8oROsuHjho1SNy17VcQ3ms4h9/hgGBVQQ9jC
+lYvSO/wsIWnphCOiI55F7pgYJKSNdVX4+UnHXrDYjZtky0bBwrwNabAfeFPqD7hiErwgzJEXarb
V9tUylmC0gBra0cqMmqNdLmrG68xO2uOPyYJGgY51MfxCEGpBoAORd12rLszmi4bO7Tng/ag3mxG
EyRkpv+gEyffEmPyEboAS9avEY0eTf7SO/peRzm4xgaQqdfHjfSPG8oUqtMgATg8LdCVW3fEkOZg
CWONBeej1DQg55Kjh02d6+ABDDT+L6wyNUFoC4KPrzukPuOamdk0oHngmCu3KetJMt/dLtMv5EXZ
o2QEtWim1/l88UlYKJL7qAV0Ghr/+K3IMm0BJPAp4jyw6GhTI0mlhJeRwN5wfxbsKr6ew6oo47ok
8U3fSyiGZw8dywC4o0mFW7kekcJmaMgheJtGOP4TNVxZdVe0Jc3OcJTx6e8aVDi3GzKmZJL1Fzc6
muXIRl7f/KIeeVV4Icedwvh59t6qBSGrhnGAt3YWNR15aK91bqWBJRwemctqCCUjuo4XzHEFWp+t
BXi6WDtR37Usx7btFCFKeoSEyS4mLlvTcdFKozBuWQ44F0vy55twL0MAcodtyYHn86CFPQacp0Qr
quRoWbacdz9pNw10OKZkl76wE0l4/E+o0Hc7qY7kTcgvjINUTZT1nBEznl++4JFcFnUjHOa0id57
HO5tVd00Ct+2tFB748OqVJ/DJWZ2ppV0RvhtS6ld83D2+4jnndOTjm6rxpqczoONSzeRcUAqLXyE
5GvuybJzwOUVaoKvtA24rfC3kjvZNBJgRDp1plypQRE7fol4+6XkH+R4WfcxbGTnE+U+f04wqNEQ
EYLIx9C3sVpSELi74IS1deDKzkflZbR5es2LHRUApWjGeXO42gNSMS/hbsZNCbC/3ubTqxKKzs6r
68CVSvRFj02dMBz9wEhxyAOwa7LOvrObOH+io7GYQu1Os/0CICiYAzIyq3r/skAtbntysIw/6J0m
PZ+7sjHoXvY1zeUpHBTaul9lOKC0KFQcy+m95u9Ry1DRP9Q46TvwKYcmDU/iVvTtxWcHYv/XmtFD
EGwTKIr3Z2J+ipLEUxA0nV1vKV9uuvfuBWqmykTW9WS811IlZajGguj9h6H9PJ49B3vCqpuNCjga
9fdj/4Z6/YZ+7GKmmw77I//Pb8E4GtjsIHFNDg+CYg52N5Btq1FKGBapQojmmLL6oq1uC2MRBUQn
cQ8P/yJZASsYeKF/2wwIAEpi5Qre3UjTsGBB0YR05tbzla6LjnbLjjchNBi8/8sad3o24RLMRDtJ
Vy9m2m80gduylU4yihz8QWQbXBBA088ipJzreaWCzS8wzAFSP8XUWPw+KJ2jS53UuKlkekwnoF8O
JJBnv1YKICjirm32yrdVMG+BM2j/VpyY02xHuITklFoRMmhcrfGAkz0+lqNxnfuA7tuxFZnV+RuG
WvUOXrIgi23GuigeZiPAzcNl0DCJsRxadiuPgFCd9we2errz3fM7KeSzdYykx6CtuNbRpa6J9QRY
XRSMBL45MAvI1+QCpBZcieBSKEtNtJtC/JZKHLSyZI+ezQKrIy44qSKTpf1/ocADy9LGodNwEwKx
ZOe/tLjjVA2tyVw8v+371UMxXf3S+yiHYYUHcSLeERycfgJQowi5/iZu7B7xpBFDfFpcbtf04zFr
E7wWMb6OvFQpjniiX1r3G89LIVptINA14ZFpgCnItjnCjTBW+T5vTKgN7enMlZeuEhZa/xeXgwXL
0NDa7QC+RPh80JA7NTYn+TmvYpWolu7Ah0VdqaxHywWKb1IyjIbFCIf0NFuAHGPVqubR1TtBA9Vq
1hMXY+39q67maUC2YxlKzxBaTRxtCh7uMnbtiD+epWboOjU3ILlBhLl4E1t+n64DnCTSOzoy4M97
tfR4KE0neVdiynRIrwm2Z2tDunWDFKBjA7PfHnoMzqIBVDuXX/3vZLJWu8ZYPsiOehjMZfmK0qHC
wzOysa+zS7ZzkKQxOqPTgT32jpQobGSgs3U01SstexKSNVJBcS+C6K7JpHKJxIAuHOro8+yFEW3J
Y1XOldsuEbko53Iju8Oc/0hqB9BXhXugn6mY0SxshRBZlfndatrfcrhFZAoahjZnztrFPG4ktlGd
yaG+lIbQcPC/hVZ/UcSVJcac1NIEEaAC9VcApOYf3u34kn7O0vhsBkCYePb5tVeXevDh24DgV8l+
NNHEPJWrAemIgTLKNpCzrVk2aUd0uGelAKb2I0ZSga5L4BSq4QE7nYpTlsAqMC8SFXraXYKs2wXU
hgxqDPl0e2FlY1MXDHXrOaCIgUBgbUIC6en2AY0lytNaJRqL8t3I6O9vtPh93nPQ9IMid3U5hJ4y
Os9YaUhJQEbMBBt+lBmxtG5fE/PjY7fIWTg7SHkaq1xDIE6EEvGGiJitqpBE+FcDbvwzbSHpafp7
TmoChXRYvXbAhk9/3NrrW/ZP/UaDValb/WitqoGk7QDjItrpiRsNBwLNFoyylJDxBvN4WZhPDO1i
eifxJ7Xw8aSkmAsjyFByZQNxPpKpqUnrLijAGGWDUSym3/IgvfxHvMm+otW8scsBUmVMAKSJCpEc
72FkS/ofqaXKEIz27rxsjqRb5hi1+JME2rSeJ+m6Z0G3z+R6HSNydB237aQdGG/Pbb/MZvfHRBNJ
C/GFdgKudznwMgfo9SWXzJVvrNwPkWSjyplxZf5yOO0Gwz0u+4YYgM2MwYHsyOnpHfkBAK2RdGgO
ZgsT4wCoDvrP0bhU+pNC9g9n5iOkhWeWs9yFa+gppQcptHwkNy6vOMJLc5eu6Qc3aZmmZihlPLtG
0Et3nnhpFaUT2PrAHLT1pDlnTFns2+AEq7CWovLOl8vLTX1xn4OTBn4ZlBzAdFV/nc/1Fnf/aKrb
7ITJkkMko4LV8OrW97u+ZWDx3m6ZcLuVU8v11SPkhPf0SX9alT98a3KPD+OKeu1JBomWxf1ei/IK
o9sOPJDI4tNBCMhUgIeMakutbt/ih/z7/sChaexw7dqorYRcNPmfytVLInEpPkfd5BxhAGbpsvzM
55bdSwh5jiQAZIGyZvjm4FpGxjJQ6zxilfzaFUhvAxTDxUnlHBhapd0PZeNuEGb/y+TdDx2zPdXM
gTRFUXy6YGDD7nAUb/pcQ7tiXXzwoydOwbeql4UmvBOWH+iME/EE7Hn4y/He5xUK2xPTw0jLpuA2
DvanLXqs/Vl9gKH/KYiQ95geYFlKDdbIaQOgis9REv3Ga7o6E6ft2UlDPf6lm5er3+m3vc4UN+pv
6OuQOCSu/+PbzbSzpsGL6elGW6GEyM8FSjgc29o6Eg2VeTLtwShaNNmrPR8QnD4fc2qzFIm5mAUS
+E7D6r5S9y28npRX71FYkNU8JUz6LXji4GfUoOYvxwadwbcFqaTWPVrfIVBBFCICiFj1ApQA5um4
+z0lob8MyUPhKnGSwT3+gQn/r2aCT5FXW4VIuBH8rVBMCDI6ZOP9+Q+boF2Ye/TzFTCzoQRr3ris
3pGufdiVveIWy1f9dn7i9jP8fmnm9z2v+3z/eCloLyJWkMQvjad+gMEctCNm855JXQ9J7CfGB6qV
olyiVP02I2qrAlmPCsGUi2PUaOjm8eA9na9CQvH7k7GARP2BULWD8H8aRE9L1NsNSTk7W+lvTMnC
CHXZb62s0QEnwgRpg+mGtSXIyuKuqK6RTII0w060dzoS4h4c0GBa8e7Ag2EqgfSX9LAdfkTCOe0K
JTdZChtlto88oDNejbRtYMWaBa6k0GTfZulKsakOwmkfmeyurv0+I8/DjWuyKvqP5V7sIiTMJN67
3HSmePMk2IeQvrkaFiu31wfNKvfu79BBdtzvzGtNGMZRham8h0COzv2+eWceKoBLWe1H7T8utBg3
eIA3JlJBSBhNpXespmHrv7b2e9qYZVLAO6klBBWCEmk4XPrlrQmrspfUrPTLSKRVq/zv7I7Mr1YJ
+11ut/ZX3xy6ymu4dFwvs8e1EH1oePvGyhhjaP6+Ke28p13rh7XTWaFMdfFK0/5GoIMDjQDX5JJV
H6/IOlpw0A9xc7OnlA5qfSUqPLXR607Pv4UTRPyZe6aSV1JfZzl//sx9S8YeT+0/JPu5TGS5LGso
vnf+ReIpFcvvgSvsK6ryJ+im01AZH37O5pVXBKjFJzT83b83QW0KvTRoKWEtLVH72AdM4O/MWp/p
FUv110UG2lrjn4bBVW6YQiKELCZikhgzwfNpGmjOvx5jo6FANJHbXhlhtcns7/EK5OsExXYA1pGm
FR1/MYu51bVE+vjqc36kyolN82iN6DGn0jqZ2lxZByogk1z/daKryGaitYr24Av7E8mY++WZ+Xn+
4t0Mip4U3FVUR++/srClE2vf7GYP4JkXeGPV2FlUli2LXNKCL74WlaeMWA1Ef6jtG71lC3fe7c5n
5GJ2Z8vK29d5bpq8PJioC8Gz+ewe4RIobjZRGxcwjYnZVtLVHkOdaZ0pJ1Myo4312DxC6RFUlqxh
3mOd7dHJz05QFNJ68MSYstHqpx7KclyDzziArsorjbhHo7XOV/3ubXKcLTumWhV1vIBwYQo49BZt
iF5uVF++DGrdYJ1pyueVjkC4uYbieF1XVmcRN374kLLkmA+WLgJTzHt6qv6nfbct6/rtuW2uzfiP
0f1UMZt4lupauOBGJw81EeiPl1NvqF5eOF8yrF71i7yEJzdT6fY18bjgoClgeAMAFNDoO1ZNyjf6
2+xkTB+1Vgj13yBU3AVSCykQeYx9Fhv3qTgz+Y8kRjloZkMvMWKA56zttE0E1w/fz0EpdXuta43v
FIIQ39yfAqAllvgWUGIbngOo2uATyNioi+OiHZoQ7MCHhuFkLmNmZ81bpi1ATOchm4y4LZz2zmoW
t01enN9b+E2vO3IW/IqmkYqnse3Tp1Uaf7BgYE4HspFtwrhPVOev/98DTcuCu5PezHwZcvSLHO/J
HBv33vTetmD9ZH4UpDAULHNsNv572xUVki2vSjDSSZzachnRzOm1SQRXncn3IOPcSQVSfMWd6XLe
gMFxRkz9F8ttOabuImjLPwfNBtcG/+moTMIqIID4ZiFGUmAuYvQ6PbFfinzjHag2wPrYovQcoKR9
VH+YkulZ82p4XcBy/ohxl8p8Tk/8FQ6ITJvQbLReAAgmZdRmYfmAL5IF3ApjpZNeA27hdAh4v9Pt
iVb8NezjzspTBkSniGHf049UgcT44z6uCs22420JDxfn7Cr/uuMK3FDaZDUzUf9mVtGtbqctjibJ
+WNpRW9xsf1m7iaR0/WVbtpnpHAnkCIqE8kUUFolrGA8j2GDAa9Lg0MB2lXwJc8LzLfwAORKxmXB
5AR3KTOYGY8UuZceApgFIAyY7skNCdZ1pSnE7lo9+mhfW7Rf56PGzce/4V6nAOijmlMMUuybU4Xk
87VuCFSfscEXnkiuH/HMmFpJxKsgSFhtfR2SDPmG5DGJNVCZFes2aI1V48TsgtfCRxSFcLJjNHJl
wJm0xkBF0vl6ttPK3D8r5nZBhJmFI1REmLY0Gft0gFCdkhnCBEXiezvlyiHg+qcGA2MqNVyrbbf5
ojxS22xYV4ixbVbEIuvejtV5PNZy5NKf/n26j+5vxo6Wv4YAXp4BmQ4biYMyoiB8zCW041ZnHNN5
hs2zZDd0IoDaiyqKXyc+0bIDF/3GxiFjMW2S5RfqGLP9ENVBgZURBVwziUvqrbFlQBLUfetSjLeV
nGpga9RcKRDp+QYWlUId+Yef9M3yP69nQ9WvTkvemmqXvhP8hG0M6DwHWB4JS67Kq7KrFapx2I08
e3viDMHIOqIBW5J3ywAacEYeAySf8bqScu1RX2yb183jhJeil2G+/5zY6AtjiHuSVEflkWhOxTtk
tYjQv8jwtsJDdNAV9JTHIOiDb0ys7MqW4lyxOpOK0bM9BthBiSJWZ0odopBnjgwJaKJjSgKDzsBd
NC250XiNG4+gbnmmDV82RREuLlXhFrGGvXBRbZkIbOWSXfehL+AaD6u6NsvHXSe02saW0dPihQxi
PIasm0zqrAlV64SCONd4kA/yhnWVZn/o8NiFNUFuy8mYSYKsp4BnXgkKIkrTOYwyf3BHjw9EtMIK
9HKWL+yxvslc1hdBkW05FqKE2Lrx7khemui2Q3td731eQFlRuadQ75CkaWU870/CAroAtddgTeTC
VaHou79ovewgVOcCHtEHFOH6oEqR+GOV+I/hWCFIlrx3wvG+b1CW+VfWcqcPNCCRFg+UNS3kIgiN
i3koZ9KyPzCXhWnjCEaDG/JnCYn/HKUv7A1J869ThwSo15lkWLcA1MTB18pQnVE/RimsSDWxgr5R
oeuKxNklv7c0nlbp0HuKazp9CU5paYt3IoVFBmsyK3EwTAL33POzGBBhq3M140k5mokkB2isX1h7
krRfihWqKBi2Eq9ZgKmkzBfIlRgxKWfYPnN2/zrnYTfXWdDFxRcw1Ba4sA1uvfSPgv+AEqPRoBli
ybdEbGUC+/KMNXlUX+QOHGzxiyK6tARAo6pOKorWILGNOimeE9oYcVB1iDm1zKh3TKcox1rFEot8
JTBOb/ZdY1kFpWv9u70Hjv74tgNzhV5Ec7GWsPcNTpWwQ0nx9GxJQsTD2wyg5fN6AV7HyYpmprtK
oeApCHr4FgC5Y9Vj+qyYwM0RTNNDaXYX5c+ybZ8FXONEnH6wiRTMMUQR+zv+805lzftNiDpY2kvH
N/LR5aZIRRhAwzKAzds1Ph3ajlV1XAChEW62tli1hU2NJ7o5yoMyrjOb8G99a/wt0IpUopyoOZIt
tToZh5ckizblRRxPd4ymwCm+R9eSL1KmF36cHm/N8KQ74mtLpwWoLCjOMnulPSd/aU/muxX/qe3S
RpKthw5j9g7UHGW15pSLACL1gG8rIzjCSAm2xcBqbu6qqu5kv3lfPWsNLBFZc9wEg4CS6hV615UQ
NXbn6kySS/n6N6zQdByyaP2tTyL5+KlLJ+oL2tzPZikmg75OlDcQXRJef5ZmWXIHsiFqesylYeW2
/xEUOXDbRQiM9E7up5fvO9cdRLiKY98JZ8Gq08xQIyk12QvHV1n8UmkZ5wtm+4cOOEREQ0THwTbX
qU3LsQIzVDKMPX4pqYVbg0O7yxAulouUblJwJcSIS3/pUdzgoTmWLBP5NG+o9Xf9ApZ3f5hpVHVN
jKhkckBNFCBv8llEYMUAgDssqfVUsXbG/mdDl+msHcynHjYQMo+zVK1cwqM2R6v8EzRZ/PrL00z5
D8W70YlM7y8Lx8crn7HytmuaDXtT4H1x1PKDAqVjVe435f7Q0uNlE7J8zyGxU8qlThSa6jLkuX78
l34p55vCDlnzwhNyARH3FSrk1knfX8uynl1lHLTSEfRBcBsmyE1XNoRyc5J1s6kSvejT+ZncGzpp
UDEGzZe5xAoOWmNiAhNIP5BUQVGFjEbYfFw4j14Yxk6ltHTdCyAZdAOW5vvqnfj6X5KvxgxU7zk4
6gNfUhnZod8SQKhKvNxoKWdu85LnD6S3bKqSWUZkF4StyK8BBx8R8Fk5A3hgE2cgzugeTEaKciAt
b0WVZERSZsu3tsf9xB3VG5GOtFjlqlg1tbPFJx7ONYkYpbqzpbFAWf4RNUHTiso8qsUFOKqO6tJr
MYxzBUHKdpZMtt8ZT+boTUzymAwSrskIQHR++N2r8BjV4faJRiusXFbLi8qxFOPVL0ER9Ego3P7V
+D2Nn+4ToZRkycbvg61yDce/jPyGLRhegrRSMkcMefn7MYTqD9Z5X1C03k2FvAi3X7RuOyW/1nyZ
LMQy33OZyy3xXvFFG1ILMgCj5NgtqZh2G/PhpYo29obOtKn0DPLNcojmxeBG9wjwLhoR9I5V4kQ3
keIoTMno3MOxnMujJxmr4gg0pdAz3gnQ9WPjesWzuRQxRqz9TI+ivxwe+rheXIWMUr6z6rBNXrMc
A0DbqsFEHqfQp731aJo1NML/JNnO6PswSXPo8XBJLspGXdlpPtQv+wPZQY9ahmuI0cz0lBEK1bv3
p/POz+DrFtQLzsDLDNr7kcBrJ8ToIr6w0ngadOV6LXv8sN7iwADoL7McTz6v86V04/gyye88x0jo
rsoPfpohKwedSpRTZzxCUC3ekvPy80WO6umLD8F3ndl/GsUGzVFaP+cgZczbao28I6hmw7cg767D
NR6yVnELvsladY1uiPATsSCDl0tzKZqLjzr01iI+7gkugE2Y8D5u2bvlnI8e4cczDN+VJvdKIBmW
Rh4enkJHzw+i+ZeYTD9hpxDhYkG8NlwsCSsL2KTXwuP0rmYpMA6NCllfvM/KAmGRS8iuBOBb5m/Q
7vJ1uz2PxNnw1HdCSwQQwKzjinxgphF1M3H/Zq85pB7GJlDHX7DKg3wY/EOtUGrmqmovv+53Y0sA
3Q/1cV+Cq8NmINR/W008Sk9luYL0wDwbvYatypWtHMxLRk8rnuXII863yncNgEtwY/+6DXOobGQi
AzyXV7RAzwP/t1FyBiYs2gyBYoutB1Jbdq5m/Ik/dkbhBPI9VGg53s5HfUGD4Zd561kS/qxMvkqB
cOIc99DHlCy/pfDZm/RPFd5iP8EO6xHkAIBe3b3/FgwPmn+psaNoWIhjsapwXzsQdnlkhntJxmAo
f6+IyU0YpQp1qptF9+Owfglo/8DKp5wGhS7mJBjUdFHA9m3wLvwde9uajoXq6Sqnr2PBbrguIw/6
6qC5a7k7QqPiW6G6ferOaASX8w9DsPmIG+s7ncGGkkFOUh36tdN4aNUF0UhTH0AUoOvRir+esLVI
eHSPVnbiIwyeclkbfoghWkA+sryrJbLNCB+gaei+63adorZ3O2kz9jKbhwQZGTEuchSu9mwQ6l++
4l8cN+7LB2mJ2QPAthdaap3r/OsrZzLVj4RmlV0g//H1QzeRf+hkMiX1v+dsVpLLoQPIu5B2+iyJ
0bUAcf+7fQdx88RSfSzCjgbovq22tvc3yJ4JZLJlmtbFA1coDbjoFjSYLI+lZS1NPOM0oEcEvCjU
iZlvlsIrAVMrprOBRp7A/RV8RgbYwfEo2KIR+w7oOoifOMSAd/o5ZocKdm22jMdAZxD34vTXDkrb
e4QM28PJwe0uc3SNzidJYdO5N8qhbEjZZ/7coqyv78T/7e+cp12TB1dEBnNAcL5ziVDF8e1PxQL0
6u8WbOhDFJrur/a/+oNDcFcyVhRfrTb1s5DgeyECg3y6+PysX9cTLoWX7DI4Ic5xQk8TXDVEp0Mq
3lsz5OrQq6PgV5N5C5jZ884FFX3YQzjc80+BKrqPscpFQWzssh2qXPfFwYD326sz1XxG4qRNNNzA
VG5Li8le4hBBrFB6Gs/gI7uAFwa75Xn6sEaWNqfBr5Vu+J7cpBspAsZdDteMus7AW7OIP72xbijE
1dPzNQ/jvJByQWhqE2/+YqFul0iBuWqe2Aey3kNvLpKsDfHF1XXNgLHgHDXpjwMA2RbN8KhrKK9b
ygQ5A1qBS2Fxcao/GAKQqm/D+Eb532V4SqBTVax3hs93xf2eJUnXaP1P18e37K1NkwIK7lFhgiWI
QimC11hmtXNv2sDYkOM4a9pQt/R7wMl5jy2Ez+5h8SINuwUERxtITPM/CLEUaa4+kDqIUGC8x64W
toS+RrW/PIf6ZZ+cDlqLvMWppNXDSx9wtGHHnAeCPP6iqi3atSr4ygH41cf9nWcZn8P2PyiwCDB1
D3/+GGnVFWY54JglIZ/KFz9sdzRmf7DMlQwgptCe9Vf7dXervAgBhVT2TwkNeExhLrwrIfLb/wb1
1SOZTOQqqSaC+VAWp/1rvX4iMyuuekvWpzgTVA2WqjC6Z+MincYmaoFHiP89S3QjmG7pkV1ytFlI
wDld4Ntu/cvx2r6uXrS8u98G/fSIHeLqk0y346vOVEVmtqkP+u8MMjIWvL1Q2voVMZs/WVEMHah3
XMuzQ4Tsrtfty24OGyY1S4ZTIrtIuR1C8C+8jXdGKE2rPGFwKomJoV7A1kuyf6axXJL+r367WgnE
CoJHQ69BrKT73D7oKmNZN8s5gV0nh29jXecU5IDVH4Dq+w1lpyGFe7Fn9AlKXr1F06hBWmmwawRC
4j/lHDfNQOJWSDgX/FcdD1PFOgGL6Iit60Owjfb2RAlopByMPr1byaie/nMn/m6515wkQ+KJxWQw
l+dRVrPVr+tomV5Q6kPkDwc8v2ViwHt1h+85pmltsfkESR+GZcYpavN/92oZWHbQIC7lEEEJVmu4
gi/3wQdlW8x63jvzIQ9slag8jgPheVRD7tWdHNxFKc/8FQO8FJIgsYvWXRQ9664X0MyV6ymSeVKU
jEt5/GJPn7pqq1QTbKXzDP4ospH5x4JFQ+HrX52riuwnnuSfIbbaRGIQmGzkhGBqFGPUn49il9rJ
whJkRLXsL2neGOP5kGISQx5YroXD+LhaRE2z7tJo6seGeeXw0oNDDh3s/DC95u/x6wM/Ky/eb0Hm
cQO7o2fqIdfIoPHclk6xS2SgWv5Q3RnwbBU6+AO9ulNyMHWfWRJzLrtS4HioihS9yHg2QUQng6DO
mlyOgVf7kTLCaSchG5msnxGu4FZNI9QPittD9dF2UKac/GEKY305oxfZJyepBq+BX53d5fhd+nwn
oJ6yssxSbp3BE9CPBLCsVolOGd1IIwLZ0w9hUnYZLBGKFwYMqLfGfJr89NubH1qg2SHbsoB8mEyw
SqcC+ZvZJwvyyXtataevjgjoDQgOhCcTENA5s0TTEO/tFnyxhkDWNenqBkuStoSiiuwYJRPGOMtA
GSZFL1BSjzv3dEFE7o0RGaD5sa1QBLg2A6XxLBEvEzrOnFAv1wgNmQ36TdcPBGtvAGs8oPEeKYnw
51iHisbNoiKbOOVg+BR6PUoZFVg3YZUuXdHQr/DMKLnJfmkP+FC2iTRg+b6wmLlNEgxOWJ8vGT8L
2yJX/7OPP1b1ym2EHFMYTiO1/ZuzePUeT69PFWAE/JSBE8zvSS2BauPAMblLdhnldkiZKDBddpCd
akWVnbjoGZtV8Ve/BeM7a4vfJVB1DxPSOr+oy6st3IXyNbjjxqvVKUdn+2xJfYRJbEs6y+f4Vl6c
sQxM3QuGq/hVEP12W74Py1XPFifqwpfagpC48ZxoXfyiPXlzG+lWSc5wI0lgz/WWMaP/PPR6nd1i
q44t+a5Bs0cK7V+8nH4snZFDFhlresNx+Tcy0iZkhrwkoje5lfV+UuyBT28Zv5X1BK8zJlch6Ctv
wQGnAMCP4QQVhkj1KjGCmTqAoP7ii26ZD72nAIN/HlO7z5EA9Hw4rfKexusyakZoq6fCsq8f4E8E
hE7vFcpAhM8M+DSvdUwllD8IkWjD17QTcEDUdRTTod2Q7Ot7qLTrBkmTfBdDOq8T+ICZCeLZhMRa
zPoUf2iZ+YwMVDiwxXRa78V2lBMHvKrqD8wQtvv1427TupoXWL1iLuVn4ZFvY3o84+me1JoZHivB
O0T0wqJTtn/ylCEnjQOy4JbttueHyTPD03MPuN93UennYjhnUmegZleUGQivWLHDgLz37HzRFID9
LwOXmCMaAyWs2rV1tSGVkhhewvcN4uDp5uBUrx8QvNHbF0kgawf1lL0pRe4nx8PvvMbFZIw9OWoD
iOiTMoLLM0btedxGN2lm9Xr1ip5Y68CPutIFF7fK3Gf+4L12QdVynB5SNhubOxlfa9z7ExUJbZgi
JdP9zVnZmuc6Fwnvme39HqjHU+hRzPz7cGdmcFSXogcEBPQG5xL6j8ZMwOQuinpd3FmIpsvnIMbK
53L8bReLRp76NhrUTRy7SIJccp8VabODyy8+RlsF63o+XkLnYUktx8GcY/qEMItcYEDRVW6AmfcN
tPX4/NX/b9TZHa5Uy8m+IgBBzwHxxFEWRuzijVfTKiq++YurS9EfN1Pu5q1z3VGWZCAS9//lVJcP
8iNkJlXJFpCZ8TxSsvc0d5eNm6UK3QrNNkE8WPcNdDx1QC7EjDoXlWtzqn0igYsJilR/kYPLPNNu
tfwvHbL1YMX5TAFukghR6hCI7CCVa3C/fxicLcB5KkgmsHfh72T8qbuQpy/DJ1cEQpCkAEqwRVNw
62l9L9OljlZFA/Q+z1739bEuwFg+GGntejreSGmFZ9thmpISTFoqcCxhDY8lwkPJ3HDmImTVdMHv
mD4BZYY53TPHngEd/TmWwhA1qnhJZ+oz3U3cGc5wd3uGrt9W3RB2SpuroPfYNG2VU3ZisyDceugp
0ot7wQTZzDx4bl8Dhw36gyQDTWhzhh/6wUGjkK5/+XdviiVNHnP4DgBkccbQ9aJuy5JT7aZn0Pok
tfIS6xBcM0+mngrrV5M11KhTmwGn6UP/K5hXv2CCdpcThX+pJvB+N0d8AaGlrSepj9ycQUaCBV6c
CHvDmD4Wq5djdXTCCD361WlZ3j5i2e16F3j/xyivZEPex64Gmr6xe5oRxS/NXXooFEJf2uocQXoo
DxK5Djy2iMaShXHpTzvak4d7fDbIWddWHzDOVfYWTkELPzcNRdZPuMEutZrBZ+aHz7ANSlkIi2gr
8OKyJhlg5RNjqmV2JezlZetHIwBvNpoxsouvVBMVnX0+KlKmvKgj6TYIPW0fPezs8zSVTmKkltVD
neyAWLlXsgYRxWjr6Zp4Ro7Dmur8c4giqdtq4ZCNFa9IOl+v8AVGUI578SIrngBqfwU+ajLMrXvW
HtqNeX1UVX0EKFvoFuq3ZCc2QCdT6Tux4JKJItVjGzVAqE0+Vc7cg+8i9YJ06DpEA11pz7fCug1i
BqRTkcFad7pWfErCxdHll5TKNet2BTugu96rTpxtg0ZOcU1AI64IrLWQA3Io8E/DzIIRWjXd4RMg
YPO+M2aBAeT5oFecBMycchTroYtDHny7D15gEu9rIgCmJfrRecJJe5IEfNsMbyKscpv7uk2ISXvD
bJqcRoDfsWVRX26qXNNZiMTNjCoqXzTAzIpX5KKwHaN8XNYoGBtZ+5aq/aUvD3HfugoNHbOTyEd0
OXM8BoMdfm2eoxqYnuOT0DDAeUt0yCH2VMmKvPz0do40rAIcI2Nxs9USMM9ZptHAEHDfXM/b6Vc9
4hzxLjSH4zFBD+R56AFoamKvq2v6gCd579CJoCpjPwJuLHHPQhUY+9KIMJTHA9QLkEu4k+9LGCIX
nrYN2IaRCVcJjBQMkZtHMmqFMxZlh8rFR86XPekcJUk3U/rqlCbNIr135oap9IRRyNxDOzkh41Vl
4jRqlg8w375FZI7U0CKhgoosHN2ous8oqfbpsa40ash3C4pG/3c5IqeDXGWI1ki9srIY4ppBYdns
g5po1aIsDJT0mp55A/Kgiyw7Cm6IbD3G+VkCAs99dfOzjqtBwZxP9Ph3BHc5WcT6mi7tPZpclgcU
OTH3HiorR0gJaZXwFb1jP9FJupwndOEgnEHNZ4ioJXG96c23/AEQtvAAlLpql4wEUIBbwUMdkqae
ZJq5SYExXcECgzBmcSPMpX751lIpXR7VxXFTom1lGmUrCGaekQKOkUq1VvMskoipGwTm39ttQGz9
s3ZssizKIyI3Y91UAPT371UggDiyfhsizVoaEeC7V1rJlr3dtMunIIAiPbVwFvCbLpzqp3/UEOfu
q1D5RcJfjwxkVkduGZgZSukUgnshhVarS9iVOgpxRGq0nJMyopwooB+a37rW4zRwNiR+bKIkhee+
cU5G/rBu94I3nzLqgWgwwP3Vr8LNlZQFhGQRC90e4Di2aFMHpIJ2ypA+zeoLMUgCAqzBOxJGI+/E
Tw/bdj+jN3tJnfUss9AyOBcJfSfE2p18WABjN63CY/wFc+GKy7afwtLSOEGWcWGVImtxqCM1Cugi
3tXnO/Ga9B6KK8p4ERqvdDr8OMAsbMVxgZKPpCHY+Or9PGOTV7da6nfJwl9t86hrXQFAtVzs/EQ7
T+1orHn5cKM+PUmgKZybPN0LGQ/yldUGBT8ZIwNDts3S14GXuW0f5lSW1bp3RL5OujQxg25fYPcZ
BzAGRc3x5KIHQ0tT2WGOWGSWyeZXCHvxpkNW/Q2zFCosIrQdRkbbFRLYI2Summdavy8Ksw3jVIPk
AEDmW5uOk3CMf3IjWwdXwgWb6y3nfgf2F6H/vAPgAJ5BP9dZ2yljRv0xdwKoS55AkuEKBZY+nLEG
fdbgXjP6URmshaMMWeFLpyrX7xUGbOGTe3KqI852rw6zqcfqdx8IDiYhYToE6WIW4dJT+ayBmaux
nP9bMf4qOOaz9qsnUBW683OAYxouXMP+aBanUdBjA4rHNWCvjez+MsTmYvyv7MEpHm16YlKD0By0
RxhDXC5tTAac8jZo1lvjS5JllH85gRGUj2Ncc1YHSLaVtJrp3QcutcfAl3NL3EB1q/bVIV2bG+vl
V6n0KJ77SMGmJDT9wF1oBzmFpGCLW8y/+N2Us7kfvFhmKdaicLFuiqClfkDJLezyWu6RRi2NADgj
V3dTb3fZX7H1Ofknih89/rw7uPxthc8yCfnRI5ejl96xyFTOyF2huehsl0IGmQ+XRX7nvDxH/Z86
Lb5YQamKHW3gGVM2ig91V7r5Ywm4R42n2rTUUuuVrOSTf9atNUgkM6D0sWoO09pfpcldPaj18FQc
vXtdg52B1YoOAr/EnYaOMw9O3fGoF3feHcC0QzbdtoBP3AbZz3O779s6hfhbdVX/xaGaAvkUb2z4
hA/VFOuowPkPDUCE/9Zsd3rIz+wWwXMJH0m+ZqH2dvzisqF9af6afffVJlqI30lmK0LWADL9476v
neyvlJ4VLVMm+J45pbU7yp28gIGiBb/lBLYapokk7MrlBJzSSU7FU6RJGNSXRuzsIKvmpKtrmNh7
gIyWeVJhE2BwqbuCrEdl5Eok1r0wGaegrXDQthY0oZbAeu4Eci1zGmFqheka7TxjoFOU41eDTLon
6gQB75FykNa04jbl9eUkZ8CF626rNUS3wp69f4pwgRrfley+ccfWSN6J+6taocVdJyeKfPwQ4ObL
tSshN+lEmcH6rxQ7DQyUBkjhSOP9ePKojF8eaJ++78+RnS7G93I/P7bpETjwr6ppg9guvgnJ9AGH
zdb1oziuxxB2xSm0TM58WTNz45dqlTafu43XRqxcR5ZVKQjXO7ZoBYSoFFQ5vFlvUELOBsnEdW3k
iDtwBKhX34CDeGsdkvyRN80tCGiHlqMVrmy5py6BQ2TEK3J3zJXvppnEt24wnHz3hYdBq63zYNVY
BPA5KNnOlarxY6uGQBk40czzTNGEbRV9zukUFuz6FCZdFDCj4FozRFrAqSc0x2YiComnPXnZS8kG
YxGrQwdzHPnAdZqnXZStvVqvSP9GGTjrrVjsZINyObUk9OCFDuYd+B6XahxeV4MkjFtO3nuUsR2j
uM5EASuRE6a31pLIPaRN7whB3GNcmniijwZ/ljGfwxFnoU7NMen8+A1caVxhsAj5ZqOcWeaEiRBN
kjLG5+5Cg7G/+zqDrTZTGPNTduT4K+wEpVzhBcqYdDudOB16ewwnl+YxSL/pNt7tN+lgfy6Rj7No
0POQ/uRUqEura1KqCfi3WanRMMtg6d+hhP3iUBuZCIfryrkh37BBrLabX8MmwyPZ3KNNsgpRd8VB
OSpxcmUz7CiSaZBehFJhjYI1kU52oOvtghedIoCNGzLUHYkJ4JcqMweA0TrQjUZFMM214MLX8+xy
5x0o+2mXe86Q3T2K842Afz9MTQFNSp/O5ohdvPOnHArMDza9r96zzXEOFYSEB3GZi0MpXWFMbYtW
VDjALucf8rxn7kOdvQD8LVr1yPXWRCaQVHTtbisYUTEhkEedn1TCKGFQuICMwMXqQj/wXC1TYmGW
yzbZUngpqxVLgv92j4FJq4zzkVw6Ka21DeKL8WUIneIBtmIU3UwNezOhyng5CeEoqbtOl+jFeNkT
KrfXTtgJOwfsQWohEdSfCAN6sNHtqKSV7MG/9n2lkrGO4NTxDIgPJgS5pr/LWQQGOrnebd8ZDEHd
+VQTN9C3/Y3v7zC6Sz7nGAm8PK/HpTpP9XbFysjaRO96bCWyIsYDlyBL4uj828oclxdh1WFl1C+s
1zTyOlag/8L5PHsTYP2uqlOHgB16xax0WGdJz1hyEdtUW+7j4bnBSNs//eCC56ZrPvPVznNiIiaj
VfTUX8zEHIopMnQAfpHQJ7lRXeCsx/Qjs6Tgx0cHA22TDg4hUMBNFT6PXA4bM+L65D/f2ebugdb0
nt3CWhilLaeYgNoIEu0Hq9704emu94/4/GYIikHQ/LSFa46UAAN3Ow/CSPcNh9+unkEFyoXuf22g
56H2OiFnB3Dsy+ZzbQMerXRBF0F8LZhjudEUb8aJZo0Evl7BHoaIaD3Bstfe7ONBpb7jol3XB7n2
s75cWMzjCzFXTgJJV+Em8HVrNuwVtxm0fTM7wiq+ewSBC7hofIPdfQtAbDkmvTifMlWRYTxgQiwX
bwyYNseAp+/ZWxR3ririb4lz1kIwVbyGSYfvAjSFeh/JKo+dfIeEqTmw1c0WXriIQwXEGfzdkE56
ILA4L90I2UVQqo74027hJmLBbbq+Ho5ZU7ACofvzDGYUFhqbQ/KsNoUzPh7OofyqXxij7PK2FhTv
uRW4I6HZfNoECOWSJxt0a3RrS/B8Tp5bMHgi4eNYW9bLfoqx+3Jyhp2DTLbwu6SYXDW89MNaSEOy
bswRJ+BhvQcQuC3/ujrGKZv96LOkreSYaT0Bjwgxecseaur0A8T043/lndBKhjrihACaZFsL8pOQ
dDE1qA0qqL27nyNUrESIY9wbGxI7ERL3OAXgVKlSpr1Nhpiw3+6mZ4FjsFs8vp69sFJrzcvWusGJ
GJuT3MYSN+QBEetXbmN0IBmhVybO47J4Zlxv9uRGulUJD+dOvhQn4RJD0BmpbzK7Z82OHyJY8/dI
+z21f+T6/rWP1z4xU7QtRuk5LiTlw+SfGRoumuce5rsBtRGzrjz6Npv8ZSZeCyzg+yr5TV2wcdC2
JP2K69sEldE8qsLZoDDqOyqjjTL4Aw98xcXApuuZA1KIbv1mz4vT2a6jhfrkpRJRlw6PqvYHvWM4
X3b1o2XafKisbAIdUtQAJjl8Z6IFXOPXpYo+TXm7ubBwDsOBIINWcCz4ZcxHXjQDEG1DHdeHb3Oh
0dHUTra4ua66nAIHnyc+5m4aChvMnx+V2B7r82lUVwAu5H2erBcVThqU8CoS8Tj46C1wsZ8mhCy7
1s9WPcjm+a6OaWZC0rKSGvYOm9zqeeoOKY6b+IJu0A5Yale/TcQYbmdrFnaCNWgVXUTSZjTGGCMV
edIWxpF6TmjPaBn9z2akt+G4IsdC7WtEWyVxbTAzI1mbG8kAeQQVPj4HZB85n3I64AxB1Cajc/vC
t9rklnbTtKcuJd9r2Zk+52IBXiWNDjDLMRxDT9PrMFTmBysUBZbmIAgPgE977+NwuwGtzFMYk/mT
sgr5k/CshZkaL9FNnGKKnbiwYlv8Yi7H+hd2W4nsIV0xxNlZ0BMx9HLkKLOUgCvN9azMO8N3culQ
uJeeFJ3VF6dhUsSUzmZ4HmzeQYuycrFXwlPzOWx+JYzbGIy98IoSBKEZPg+IX9CxYoXGiJVEBEhZ
OHc1Tcn0V1wPQXuYSUBJBKk/ir/yDqa8Y0ZaBg48u31JNPN0wHgUuQ1DkAOnWfM/f89Zn/3tR4Pa
wvHc8Hf1bN2Y/ARIKiI3fLb+USxWHUB5WeQ6LEaU5be5e4JHEftpG7vAdg4FDe0DbEU0+9tubtKX
u8KuVFnZ983Qj1HbUfo7s8deKPqcXw3luAxW3Ywt2cv0MUR8+YusSZ+DOMu74By8BrLWF7zJ4K0A
aSt1xZ6iwD4qotTSr6Buj46duyBmHdsoW980JgZTriVmBHkQYkT39xJOgsV+ogDjZ6N7Jur6IUE3
cd6/eV8sWj+BKTM8YZJx3V1bQQyiSDm69irm9S0MzmNQ8z5a0N6EkRfthL+Li9fvPvolUMVRmmAl
KjXpKZGUF4hlJ+9nI0LuA8C+hGESTYDpj+k9sRp8AAMwWFYtRBAdBMPxeu5DuRyYWOINjq7YOHTp
FYjwc6JjKxPnGeAliRuVZ2uY2BsaV+ZElFJCIt6vGJQGNDP7FxfHPA3E/8kT1l+8nv/8ZN73FEnZ
LFTuI+1thbrxbK2BXlkLKbPRhiTw+EdJ8Lq/LXj9U5L9tWlZuDFHK2MZ42YgSMoYNpuASJBwQvPD
mF8IFAOGNxoc5cVGUhvlWehH3u5CwonVDZDKY6dOSzPoRw3q5Af+gbu+JWTbz7TKisw5ijVtbZFK
zblgxXmFPqVGsqZOf5UfPu9R8RQlCaCxCWXs3N6n00n5jehVhaCabweGMQvxNpkD5RsoodlOKhKt
a1o6uJD0LYDWrYiMuzVjE2uL3caOKuD0GenwmLanKswEMv8KwFNSq3JXbimU93iQIH0iDo4tWWUV
lT8yqte0GnwWN0t+ZGjo1mOKcouuGv9Ebp85l6PWmN1JZAgJlrx/XaSJg5yUfVKDets6qoTwl47P
2QSXvPBOKBi5bcjQudCBFlEJEEBLZWogQrdXViWOiu8gsH/4pY/7SlbVoW6TseUZT1QzGhuOLE12
FWy1t/UVu1yUycModvjvIeuPijAXrqGz6DyvAwrEAq8LbU0lDhzPOdaE8LrbQsKx1G/0F21vRIAB
XBpKuY7Z+xSBZpzvKI1Vsu6clnueMsv/gNTue2fhsa0YgU2+9BIJ4vtd2bZg48sS/R6KhHur5m52
o/rbsT3Iz4cPAKu4YGdvnPa4M4nM5eMHwWTud96TRh6IAmYj+PdOD9xGhdThKvmqJHX6fimcur5R
t/aZ1G5qJ24T7k3g/Cu0Li6PlUD5xr2fsGHOj4sonMaNcFHKI/9oZaO7DogQjbl+uB/leeHeRBZ8
D1X4x/3FPa+2z9H90nDWgDootAxtXWVpQccZfrfApglg7kN3VynUhhukv8vHhwVDGXtbTu11VmO0
K3eO4rF6/txW0qvNaRiH8adP4ccMBIvovP6WCnSgk7D+pUjJmJVTyiDFdpc+u1Dk1D3x4dVRkXnr
mYcC9IDtMGHCXndDtA+B28NLF2w+r1xL6OzQMEXayEsYEWPCQPEO57z3fuLLOQlmDc4MNPIlhkDz
v0Pby7BW+UvPcQNKAPdUGNf1Q4xKoOS72FU52O2zstBcEgNvFpUTQTUApavs2oaR86z2MOZoewuZ
q8pqEOVgYS5xEK2fKl6Q5ZXcYqe8eB4xOxsEgQT5KnrpgSuTtZyUvHhZfKw7RiOxPAf4KajSwpr2
jebJGFezpuiFWGCvAhvDONtc2s/IUs2ZJNxfGQVQr3Jn2W2jEygIT1aWGswWbypdiYhldqQhYoaH
0zLVaKJeHd9jrcNi5WZHWnYEFkwD51H6GFt2sRrEnEOpc9QBULpoIBLSGp/VwEwI1QHSN64OEyx5
mmk0950+X+r1itW5SVPLZpxloM+WLU0OK2DN6Q0MYwyCp/j4+QBd72Ybjdp9QJ78qKWboKCDT4r+
idRk4Zu3TrKlELGfETajL8I6cjPMYM2sveyA5ZdFdHg6jV+OZsHvgLOL1hzDCVklzLhVkl0q/2YC
yCl33+zgfVdZ/N7JAgtuKKkofgc1XvQyWfg5BdO06yjPjRK5BbLwWPU0nRDx6PiBjnwQQPx93mgV
zjP+JvhNHnCL9OIeZhjF9OaLRAW7Ctbl3au2P0QILYkTftJ2MHf5/OB1WeGQuke4D0QcrzDJtNzo
u0R+jBV2ORgMEuLRoZppC9IK9L/E8r8kdfyQP50WrgwCvXH+pMHw7jahHWkyXLBKc5Cn9WKgCKEC
3D1rU8fnZsXBCiOaucXo3uOgtsHQMB08hHu/FMOj6cZYRQyI43q8tV29sSdP15ZghdkxoyL1zYgt
+AIQv0R5srqpamRNTVLtngfECcHRJU9qb0atq81j9EZ2PGiDZXX2XzCrXlzNAjGBfJ5vX7zrrNkU
+eFOuOvPD9eslIPpp53m4RQNnVb0s5B7hwNO3hFuHMas2EWMm7VpZh04CFunkRJNCRzOUb7nc3YI
CugfNi+M79QuBT4o/jXbTuYHJ15qLSiwOGX6VpXQcRwft7PhdRf/K2n+rY+n6uiLrtGRDzmDT7e0
SAZNu8oYdyGz7p2rSD8CSPeFAx+GyUvF/0JXgRYNZCA+PQQuMjGMlezqbOCo1fev6oPIBDTFLJ/H
oXeo08ZT6C4HFKuP9sioPNQYmz3WHpS3Ldt3xjgNAju8Hlh3Xo4yuawwTLfnnb5DdXMCDh5Mpj2h
FdpTZFja03v5AAxPA+otmHTwIwjPInw3DeY/5TTXlRfICGCdydnb4Yj7msJjDi3sNKkwCMDbG/Fo
vTCBlezawQOaKuifrVNm6VdfqFI3bv+nng4XiTa7OjtU1wPZJStiXYt2HSaNs2yEWPFDkugMSmA4
67WDLTkzZDZwkMjSGJxAGxjDYgiRDzJ1FqZib4jCP+4BOd+QqcEqMlBuBEmf1888b25BhMJcqs6f
iukENGP2Jl2kX9dS+n/7Z/ZBGt3lwsYZfFpN0ZF8podVVfyiNRuC31xkwM5LFghoQS992fQETZix
SuoxwVRcMfGapEj+BzPKZJIJeEyTS+wI+GGoxNS5gkGOBqyK+Fz/KaL5l0U0WtPR+JQx/PCxcd2E
l0QhNsxIRAHguKH91hkzwon0EJLNEpV6LoHdgVIWErx8pr+kqZr9IqeBpcBqmG3FZsYBPTVbnsy0
bwGzIHFfrsFUzA/1DiaahIqzYXHN2fqBHrBdnpup7fbuEbHDUwIp0dPpVwjAHe7F23dOoFtKDDvo
NOcpTF9b0nN7E/3X4jWpFMGz11CGB5FgzgU5KIgRVB/pAHSZOcM5FNxJOgONZm1j7lAZGXILbQ/W
BTkxUMU6DLhRNCIx9U4FxKTpzAqp2SJw04I6adR1HcYcQvGUiGLSDJx15pwP1DC3DEQpeksM/yH7
qJZB3kqQDWs0PMI8D9SQ0eSWW9qm7NBBRHgzqHStrtp1tVXJFvEu8W65jcz8u9wVwW7YNHd0LmLG
b7E/HlIcxXHR3byirFnHipWIoLwsZfru7Jlt41gVAv8jGlSHe8G24T74GFY0pK+lGJDLwIM+z2MF
zzAn40v1DtwnHzb4i2feaSALK7hm05WgyY2YBRnvD+vbjYnSzrGLz8lZJwdG4HEG77uA3vvUXOto
qSmXl5l2Kq7nNi0+kOD1/haatJb/WKyFQ09XgO8em7njlrTVvPlIqjn//1Eb//xcZk1BFZs91c7E
k7ZkR3GczPh9NYKctdYlL/UrTKUdFY9Kz4mJBOeeJEYWt71+1cV/BmU5cV4Rz3KcPWBlByYnlBJW
r9nNtcAdhNHQwrzDZFrYsBC5FHgVqOsj6a4xFTNZPPdX7i+3kDa6IT1cz7vRo1vUao70Py9Re64G
YXl2oqcUZo4qqatSgdmucxvB1eDHc5rcuRyzy0a5L3j1p7MKUKTKGCwWHvA+URxYpy0rW0arxHju
ixbFz1PhJ3QVRtWgYxiy8DpTpPXiL/TgXahYqvh2uegOQ3MbkgTwk95BlTl9VPeENau3oXdJO58S
fw125mYxs3lhCaC5qyBaZSk1bDVYUJBPZ7IMYm7I2eK7svZrd7Lx57bmkcp39NEXJ0TWqnXXXs2b
Y3k+pMsfygYhUjunos2FVJuc9BCZvS/MNR3qjLFp/xjq6mz8NNPhSa/SvPRpWVxpFyJjOmASYZIo
o0x9Kp4LwKqU1QFcMKZZgsms3fEP0KF26B3C720XYYaMtiyTV76vZwgP5y7oyxOxM+TymBuSYF7S
ZiSMsTQRcsbu5prdjMvOQq4kMfcld2ATUiHWwyIwJDVTIQJ22Oz+f+xkIMEkupobQElNjBx0FV04
dqktJBjKW+ThzQBPhPWvtgcChbuzvYuqHbDHjAFWdbsyHeLY/VcOe/ZpoCeaDy9LsLmClF/qyD2s
hSb/uKDZqPY2pbe+wtd66f0kMRfZ/CtvprEFqfO/ufvn88l86IggepgEGI5G6DLllqsAa/9sKFUx
sW+bPQ79aGUGinIvfGPhGpqbCfzHjHSY1nWZlmI505AdZ7XmAmpfYr4+ESEMFes+
`protect end_protected
