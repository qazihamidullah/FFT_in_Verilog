-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
aSdP+CGtUj/ATPSJRSKhQsIUZJqPxvwRp05YhxP69gqtS9LDv0hvbuPdBH6ts8y7xLWebFTFghYu
9mNrDNrIP2Ws9+1ZE49bHXFSjztazGbHyrUCLx1Hm1JwCBI76JF/Lo52APMSIVvb7/4QaZ4Fu0Id
cT1rKz/e0M/DEgZqWhGEbHgXlZZuNpHQBodZra5XseAS9uuMoOdzDNZQ2ipL0GKZFJ9jERpCG9vz
e0R4TkLeg59bTW35Yvl+lRye8vZMSytRxyCtpPLafVkPoI7mlNrIPVUf5TdQA/ujLEcjfEx63A23
aYVOacmnwdGXjhI2e2N/m46GRYxE37jgGxHbJw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18800)
`protect data_block
LTbKufJVy0n3cR/PdDMnxTugLgFX5TYngDqMG6RFJiNtOXPSjEYLoMmTponsFG3PdoeLVAAZkR00
pd+GEmLTaCDIVp+hOLGIpDHMlGWrG3PiwdPyraRFq28NUwpo5B2EpcdcWtwLEW8+F1SO/uuAhucN
55bDODl+cyvTSwMzWRsliP3gpYkJW4mVbqsFQ+B9HQd2uydZ6xWo3eLIjHb0ZclHfCTVipGldY3X
Rbyea6YoaAuRVe4BDOotYLNbyTh+9byNN6wCdyhwbebioE1tIsl2xrHwBTl6kNULnPhrH0XouhPT
vrlbb4JV9io0JEwyW6YzoJhXOR/wfRWYYsjNyHu/vrXE+yaiGOVLHHjFRIol1CnBxtGWb38/+PoN
1Na+vfzIZTddRly6e/ffOe4cMEDHvLxbnor84LOVqgjZB1anxytgk6pZhG0bIlkydUEHnKvxpTrp
V+RrqfBd/IEJpGdrdy+i8D/wB6G2pRjwfytV6NuCV3lX6PfoUorSUSUkCuiU28SquTA2Ybf6Ezcj
H5DOFRAifvmKSPGy1TE9xFt2fQs7V6OdNXB9KAYRYzh0jqD/tGzjByri2hWkNc/hXFwy89czcj5Q
YflG/KrIu1IVOMCwvEIFII0V97qMLz1+z1aRoaB7nWyPxU13bcXG9r3L9SzkZFrtitSvcRuGpM1H
Q8j/pv5130TwE6XhTzOyHQ+ogdq+wU3vQ/aKs+JL7sSCPHTn/QAhTG7zfT78RwlGe+Gy8zlJE9Uu
Sgj9m4HNbt6x6Q9o5jNRMjlnUN6JTMBq9bMebnRi3XC5c4o3d6XHd2Ep9uG1Td0Pfw5qfYkGOvFi
m8s6egyp3gyNVc0ttZz5WEJUyAerWd6/7w+OttQq3c94CeXHKmdymQZ30mdX3Jm+gImWO9U1oqqC
5mR5xz5vZ3EW5TIoPaQlMcNY4fwe12W1TLdnW4R3RMmKg8qfc1ENMP2lvK5i37H9EHO79ofY9+5e
CON2MfR6xAdq8x6Pg4BsoYOB4Co0pi2lKK+yLukiug33Xb8bJAIgc7rLiSLkyo/FsCBSAMYa/eM6
fkeLplgK0rdaB8a6VpqQj+5Y00X4Va3j9pmnBUrP3ff4KWNVGSUE/t73c5Y6AfM5ruIvg2aYi4gf
MGwLr7GhJrJ2fgbWqppIN2/vjPYegkdAJD0jwilndFhg/HZJLN+hvS8ovKOX8PVLhV3uQA9I6yx8
Moq5SZZWowz0+fXBNW7mfEOiLOKnyKL9By4rOyQfqZATqrchxkGOhw2ukhXUyr6hEpyyGMFBe/Ku
TYP/a0LA+zV4vkO+RFiwnkO3Y2zbWmwfdcwGQhFMvTowilAKUHZbxOfJxz7Mw7EQwBMqQOSp01Ut
KtC/NK5pKor9hhXlzxSSLDwhTAoyuEqf/pRj8dPEfJWr8Dim/xhx16HojjKZoqlEYU/zYI5Q67VV
FzcSbXMez82XgncHfpvDFm17WeGEb9QWkRXnkuHHuzYt/ZhqPAoC3x9C6TKsMJ3KjN1qDXCsMSI+
CP8TukILxaQK4sD4v46e3NiMJCNZFNfsdzaf++EhAEbLayZ2EXIiK2ui+n3d9QilrEtVivON0R+b
wC5L8fGI5dsbBzx0vSexJu75PuJ2sw2CU4eZc6nzJVKmYrknpYA1wD/MhA5vn21f7E5RI/hQKVjy
ceLNCZdwnBL+cPMgevqvgVLzZkArFQxbSJfj/GCdobvjaozlsYO7nde6c6eHTxD5u/E2QMrDJXNs
xCB1flOLgedB5MJtDWhrfBHdtQptNcMRBj971e20wAX+50prEoAndMZMSjYMpNcEzmgtWZ+B6eC/
HOHQLFlGVyKm7T1p2PXD3oZy7yZRop0P+kocU8NCZJ+pqdVxorUrKcbh+Py93/mUF6vM/V3fhIBs
CK59MlpbMF45GcMwaBZOyIRIOxyII0tBMaFqShXortJaDxwh+cra0CHDlIxRuKLDr2e6EDGHwdx3
q7gmtHRfMZAtwXn11vyg44s0JK40LwEYavTC6MmTIxShVphv0DH9bFJNPHrdClrzrxzzVpPbNxJT
whpemwiV1trTPa0dE97qdrB674Rmy12/a7aCpD9O8kBFLhtR3hNk5dj/l0MON9G7hYXdh6ZbnOSM
v1T8Rc0Xhf3FxUmaSl6UE/ih0lADE8vzMBLFZ8lM4rkDQvBfYVfsJaSb8fvK2gu3kBuWWO6ESbfv
HQ3+mB7hfzTMKvBCJqFjNnNbSb15SIgLAKG8VZoaF+ulSNv2bPVlrOROqZCkvkV2rAOgmFgBm1xJ
4/Q03RuAvNL/z3nSlLrF0NnALlWnxsUHyqzWuQjyYDJQtoVcuzwOLhGzjHoq72sAkveW/Gd79kul
2IxUJwRbHH9HrCDC2Vud5j4AfRyn32P03RGutndvG+UihI4SkoLFRantb6p+c2k/jrGT085tsOkT
iFxP/Y84FcU18KufyJ9EP2WijO1t52zvNbqwFhW4Ng63CLESkKvtCxoT6++TtPc7RevpnyfhsBIQ
KxKfhCh5KScbBWJ22p1xaxJLlg6U0qdeJs8aZg+EF1Iaofu7WAl/5joslcgOQN07kzPsXwtxA+q6
O+h4iii37ycFAJNmXAuEKMKPqy1zfxd9ylRKQqZ3CSlVXSSKuA8zJihInI7YttrlaxiCowS2OZAG
rzbwBhQh4cIphJZM91QaHNs71Tb5+9Z5u8Hi7D1sletawAdZnmbOtB39BgWv1HX18PRc8yuGGQ+W
Uc7j7SEa5APVXdCj/FD/HLMEZD5H82he4v0X/BIiJ8ozvAlvuyKLoVumeeXsU11xxLa0Ly9YYJeC
QlgORbOwJ1gRGOhoYaslS3vW1SSsy03Vb+5+GHnuJBCefWBU2mJxXFHoQU02wIZVOAfcUeUrAwgG
Uo7wQInQP7VNNLosgOKfqRHxsZ61j1qMtt6KyOeQnzGOPjQrgasb5C8aghlCpw7GQriOHCnIeJTU
L0jkQxoWWiCXfjO7KNiMEVHnB7clBkzU8YThXVdG+zRDzALXoxM9eQlr1211qFucWj2t62+rEKJl
98DpFLTph70TLSxZfCguYSwOIA38G8uhH18dVgjXcXZKma8gRNQha7tQuRvx6AvLtDbu2T7beBEO
oshynqL8mODELiolM/X5Li2qwCHnDSUImeFTXgiXl2/WNgur2divNY/Qv7ypCFLkXnggJasJ30iT
Q3/i69JjU3pmwPXOgNu0rfR5K3ADy5LS+TY1WS1OT6bhyO0BlnW+trEV1m6Dp8L/RPFGVny7EHrM
bp5O4AcHrdR2Hla2sAjbFHpCD4Q+vvitn+5ytyLm/93GQdRPCSZL/kElyLwAWQto3/p4AMILADAn
oxW6RiZj0+wPTWf8zSGeQe1q/8misYKqXqNdMlrzsV4OqRUAxnOdRI5J4i0O4ZLb6zrtw3uLcO13
UuuNchTlEHYSU6VEfXD+O+McrdEoFXBnLiExEo+YfOnORpx6zPs251HGX/PPnfZgVkgXiJvYHkSa
c3Twx32qw8bB1aci+QO1ylO8m47RjUx/Lb9G2qG9TRNkZBnFAldQp8Cb9LdxUGTBC/1c5Do9SGI/
JuelTTgQi2viSgqfth/U+gUZ2+75A0F2rtc4zIvC9hP8H03Eyid7H/mm9pNRxMaJlCknFhxancIV
Y/x4UNdHcUc+jPUnyBm/3E5cTsHlJmA3AgScgSB/zK49l/iZ4Lb3rxI9lGr+RKv+CUfdI6HqfTnn
sD7LifCan9AX2Zr9GtwBP7XlSL/OwOj5mTYtZhdOgVfoZ19XPEuSqGJTcbBZTMsdzH1POf13zNTA
LkvtBDWMZUlHt3pAZrKREamV5MP62Uf0ckXNm66MbohJ9V8XqVFWZWQZUrkqywueru5fkegLK9YB
XRTCui34r2NC5GWBvmh7lhIzEdy9jSfI8LwCCqd3moxdHUUpr4DHLjV6yGeNlvdAl8ZNR+jcQsf+
YfDD6PqvKs7yFqy77vWbbK2ctAX8vypURVsbldpmwoB36uFLZg3Em9UZ/LL41uY+j8mongMKdwvZ
MbwXHtFNfRce9dJs2kz8D7dvaMq5/3ROdIMG4RpzbhlRdCWtZnFBnR3Hk34KP960Xgq8QF9qipuS
yewaLEeqVArDRo2Zpg6RMyvrYL9YufZLHnbUljUpROtAc9TIESron/B39Alpy9Q8qG/c/GZ7jqDC
qUlCA5PlNJT0XYgcyBgWVuz/YBMU/bFRdiQhwBco+Irgkgl7VfQSb+lQts9/QXIj1fx17WdxILeD
aNtPG5PoWTU1gCx16eAUYfYJqIetOpugszskHrINg3tu3dya2d/fIAhLX/6C7hJHBVQ+P9klFIIg
Ejz8xkW/xb2Wo6MvPgiUVpaEPm2khLmwZESElCzulyCQbvM1QQudz1wvODeE6/sQbtg/ZrUMMaQQ
eo+D1SdmrWlscaxbZR29Gf64naV97weP759wo8WNcS0KjHLl0HtLDnfe52uZAdVnipl4Sxw/j3Hv
iGNgYPY03CAfpFXzpKjdvPxS/dwChSclk6jHbw4tW3jevhCf7srO0UToz9zcRRbmTYrGzR02fnKW
GoFeJnKxpoZ2s5a0evjkSgYWnaUk1oQInddXR56dSBXubr6ouCS7HBuu2mCmXALRAdyFLVcyA1Po
HP9KGr7Tv5Sj3cph0ZB/5x0ru3cw3T2gHZFpMHEiKh4G0rLOJRfAU3W51djKX8V3LwNg3Fw3+zdu
+KR1YmOZbozm1jRZ/pfT6QVGlQs9K9SIaDKQfInh4mltDmRhljE5CNCuClWBmK6TNzbVaV6hZSpq
sSwMd6i+o/5gabKx7Wn6kaVZwiM+fSJya8Rn0R4ODBGdbvo2crAs5SKWOZmlzHmOazrhKZdbydBq
5lPtMf2X2RQKRjfahdKxOwmv2arWexywG8n2oLSBeSTneTgPc505gkfZBYRq7DcM8706DQf6ez1v
n8TyPsrjWUec+jRf+Nyto/tFLkXJkkb5x9pba8sxTavqe4wtfPD9izeedHR4QqOilT3i2YmvTiFa
8/q4rQH5WhirAJncmh2VY10BKwColGEQRHUNcEBY5D/tvaBsG+KChGtE7zQKH4/xS+QRZYecoCIA
JQHMjgBV1WSe5JCXdfipFJc0DCSRlAccyMu2g491rAxqzeDV1WRubfVkdAJHVXGm+cPK4V7T0qi7
XvotZC51fxyst4v6b8G361h1nXOQgVzTG7TSO0kujKhzPZRvCcYPabUTeWZ9qONTAS1K8y03bOky
OwNaZ0rJJI6zRGWqHMv/PzEShx0c1k5YNYTt0gOvnexI0rMj6HFo3NB9fZhlaC+iTSNhvzgh7Hr9
kD19cLGLAnkRz19RrCHaIfVcakhPQo6R/U5cqSdAl9AEn8XoBxDU03+fqvrhu/pWe9aaaaP4sdi1
TW/Xt3J8M9M542J4sWozhF2O10gl31Ld9vwzHy8g36r3N0WMdSu2gwOxR+adlqro/BbHs3iyxEUm
ZKeBbm3eD3w5SoZ+xq9eKEVa10cfuGKHgZFhFpeZ80A3FiSBgjnC+Q8ybE0VS06ijW0e8debSZ+d
ueSg1dVWeCzVCUKp4cBY1JHG6fJ8hzxhXmVPpbGoGaikl3tIA64jJ4X9oMK/SFDsJDj2WL3Kc86b
kxu4v4V1Y6GluvZVG4ZQPm4guCkSEc9aEGMEohfanKqw8K2HUMETlkkJ+ArHIDNXDQWg9dkbfhSB
MO8ArDyFnEUhR9mjqlvloRp7L6XwHulOnZuCGd89qq4doCBu3RRr8ApeZqEzH17T/VlMF3AGAB7S
utK0n+8fPqCqzR+hPoB4pCp9j+XyxeYWsp3yJvR7/J9oXAsYjT8sa7WFe/fU+3Ynwq2R07aaDTic
8DuaBWMywmZAfWpIl0nenpR7X0EV6DuOfo4bCXI4ZVtNdG6sMERqCJdR9sAUQphHk5FtRGJfQ8O4
bwFzbnq6IyAOr75s0ir5mJrHR92OmaLYHUsUycvyC+uYLchfY5fm0vg9zxPZo9GmMkGk7EndyqGn
IeNvFVLBAYIav2giTwJs6/rOKypJOgFd4Jh4Rm4dSiUc7hq44MxxqV0OGVN4RowInL/jGfeYybnU
bz6R5s0og4uEsBwyU0vGFlAXToHXhUVViThdcABsCktQ+qAASdSrf6BDL+wf0IsotHxHHa0oveK3
du1tjvvkQHftqWeX5kF3g6dzY+ocsMYuU601U6MXrjWsNs93srOXckIR3VSqpsE/H46mnm5vdAuz
TcV300SDSZil+FlR5mDFzBm2SEpY0+Nvn4sFzNOu7uQECYt5QJIKsg5x6Ct0YnyBUw48tmxdxoHL
Hya7/qFD8QtUYOOhqq3kuAt20DZsbSdqSEA7BDMglIkbpThqDZA3HJSSzRO8wmx3N18NTWGYfDuj
oQEpt2Vi0Z/wDOfu17/2b/w41VOZrlfTCFcS/5PAxm68/IZUEvECDDnnJBTKlNIih9rvjIwW4ciE
slNOok+9WaKuAkpYVt31wzxMsWVFBPE7kQLinBTT/XjWE2YneCl8SQtbQ3YoPvn4ncdb5F5LRhtY
d7CS/0yp9hnIwzS9IgVC9P8nHfzVB9Ct56hJdhUwIiOziBdxDFin3pJR55avgqKrinht4D7TxjHU
+F42sxE6B2QCQTRfzEPDWdBg+P00dza42Ta/VaQI4J/9dbadzUpyllfcbUz3RKnlh+6EeaiTG+EN
AbiMH3WxBdzgIw9WQQ0rLk/b68OjMInGQtNqcZHM3ttIgwRWiAhmaQPkFFO5v43siY6G623XWwHD
qWNAodIT1zGEcV5fJGz5Fj+i9JlOl4373+fSB3j1o5Te/9HP3BNFfO1bSsZWu5xENSV4YrJoekjj
PNsOV0Cl096T2wcOeMkS2EglzGI6kC9SlLfys12DQ4ScDEbMjoHx58Y7vpYP/gVMqBsIBRErnR+x
+GLUpJj2FWpB/3S07tkUVmWC1i/v4cH+NOVxFoqYmBevFgJrQxhlj3x0YdaWQrQkcs2DKaEK7T3P
Lz+NdM+EoPmCj4bvpTFdpfXepan8S3JvA4wHbMe4gjjCX0h6zkU+DO6u+4ezWElpf/PmdqFFnFxd
MD1jgsLBqwH6BcD9bibzRJ6HLHpQjo3y/7PPiKeSXad1v8F1mtZrhZ7gy7kDU4T9j4beuAXpvGfi
saVPWvASISj0M2gPfX+7vNrXqJDR257S4ppXQiJ7wS25CzHf9axzgYf7bkZdyXE7OXBGpwVZt52p
r3nhKCIKOI1GyAC/QAa6X/koskLc5vE4eKRdetBsXqFf9ysrD6jq+J6B05vPxZsduA9QRsX+ZFQF
3XF0tAq5CFQJOysqGG4/k15/pVEgePFNHHLkp2QIB/X5YeLksiWRZlX5PBJLncXFydcY1ncVk3nh
7qh/ytFVVWyux6m7FNFgKpHxMa3E2GUgNrQwzOeHRSX4AK1eDP0vMSzWuwOXEeQuyZdKYkU34OBT
CMtZNTpt/5QjgR7krO3fhOKjLU0w9lyCRcqDG7w2OYTbY+B2hV4ofmdkd7PTWOD3P56eTW2Evq4a
4c84BMjBV8+IqpQsYQdOuI8aVFxPpCiyVwcCK4BpZ5+TST7GaYT2CBwKqtYJazg+2zlAAeA/VzRx
tDnn8PxOECmRZ0S7L8fAymSwoJdwpEneSQXeTunXGRU+0pgpkmhgbiRVF2bDCbYDCcsoypjN4506
ojbXQNB3lc9jgGPB8rCvdq/bPXWxRA6nKXDlDFeA85oCQSDcny2MqSPw21CYN8sbRclUazLuKAlt
vESut1JgzrpBJtk8thpqcTnrd+lnvuEH/wVt5wOtZhM8IbDMR4iomJql93ynbFBlZWr/lFHJsnxC
YH0pmp4oQrQ9cnrOuaCNj6H3JO5+fZ9S1Jc05WK9Y7ynQ3CQ2VJW0d/JEo2RphnoU5QC5OztSaMG
KHtq77KjLC7gfteNaRCieiOXm8GKzwuPG59JvTiTsrMrQquraDK9bxFv3MydewkUqRAqNAwPkYsS
7zprLXaVxhOB9eMCIW/X0gM6X40p7GKtJ+5y6qJOLWeSDMwGgUpnfT6tYarnmxAhVstOUx/S0Suj
1RBT7sA32fjxM9TjzFuyHrka0+vB5BkDf9ma2zZPGPyUrbtbTiBo3QaRMt0BS+BUqH5lE3/1uqqc
IzqUlWSmu5SAS5X85ICIqhnszComtHp7dc/gb4+C6MKTPUxagMo+RAPOUmsbsIQYrYg7ASwNbrTQ
D3EQdDvS3C/jiNNZoApG9GdL5mVTU/IzaZYB7enwlTDn1/12K1OsbxBsF08n0fpO9SlQ25VSpbpW
/v5M0f3yUE5czubCodn6sh8W4FIDwmXQpJ7AixCa067Y0TgS9Mlyg3fX0zJPoZyAvpI64IFtnBJ6
73b2hbNuGqqjchl8tWlH+BLEkYK9JZbXKQO1xiArsLIhdlDuPkR/3fzff9eoQCN6bnMdWRSJwPKT
QCEbXzn4FXSxBtquXLWzLl1d5A6ZFR5tsUlSLi1rU1YvyKAEz/nOekDzkCY+oJbbvDug5MNzmgts
O+egu1RF5inDakXnFrU+e6zJna2BD+Kirq/1alNStPQdjCX8mPofEtg4k4l9E7v4qceaAjgzxhc/
fu5vC1d+DNBP3LXOgoxJMp/WdtMqBDawuPHtR9cl7zovjJeOpsa2CmaGZNeS/Yv8ZdGdZueWj/ok
GclffhziMaU2rWoygVTXlbrhSVVXYwy2Q7Nh60osyYQvFecVjrsW/GcMmdtOnb0T5vj7gJ47Dml7
deRxhmvTvjbFVGt2iJn/bxn5P76wboJQL5Vt38/M2M4M2NXDxTPOrKv0lwX/TM3HZOZb3vwVPEns
VL4byXfYeT/VJAaUshqbYEgtCEaemUdTNoFYU8Fiya/J4pUtMmHHzGDXUvMq6DlHHdF1XPrBktiN
SUfDDQYeEVqH1BoE075lPAbC/g8LedWztHSFyLgXqskrAgME+EcDIwChD34U58zuefHq1pZoxRvr
u06EKteo1prBsHQV6IWxavSqBSAUIMPsInr1KiIrW9NlJxsZV5oPYPIRB4y4w1J92oPM+q3t5fia
/B7/MLnuW8q0thUO3NZOOEdFdKOj2neFQpW8buzKfYJsmN0sEWEXs4IGKyR0G0XVCetsJKRdlfzH
sa06Y4bU4GVCu4Tke7js+hvE/tjX3y05+jUZbj3xwSJodeUJ420rOvLL3qrzfQneHsWdwacYy0iw
w1w93ZPymStTb5SlOM9IbJShzPLamFCxr4FcSRHJwKdu3LrBeWw1ljEe/6GN97T2E8jgYr9wZiSO
1tATyLYE2XBVoTTeVG2BkIsZSQStlncuP3U1ObObhMBCXskXk6pUQpQXaBy8CYypU+/JFPcZsz4f
zfptiCqErCi4fsKlF3fFQLsLMLl0zR6JYXcXsBFGdo0/igIUchhAZYVRz6EDk71Pkyj0Pf966XaP
FENqD0GlcIGEer6IjnhPdjJfwC1dradE4X+sgfLiSXWRi3A9VnUpjWqTGBbn3eULHGD+YbGwKZ7C
OLZNvndZx3fuR7vSAZ5oSw8iOYUp4dZOJdp1zuH6qvutu5LCE9esT1XpeBhDZlmMfz7RSAkdjkOg
9NeKdzBBKVBQ5IifwZK6RSOm6nD6IsQRuNJQl16CAGkNsJUWAUm0WSZhdldRQI1lQr8PaiRPT4Oy
9Son7EkmdKXwnY4Wd4+6iDD1/e3LhgN9Ne1p/ZMZoVmd70EacPKMllpq0i1CW50+gCCgw+nPvM6M
1cXA74estbO7B4HMFXgnCvCC1q8TH6tjj//DcjRwJKQRQTGoMO3IDR3bNI1vYYKEuFmpwrxz5yJG
Bd0EDX3lItVLqaZJQeE/fQvyVj8BnrJIQ4XuHWoCXYeMui07A22/sq0MSrYaSoUDY+NAQiphPHaf
ybPPtWoZ3ktrRJJXowInt+2pRkaMEkYOH3TtaI+Jd/KZAC64/lEUp+fOBJLvuv5h+GvPNN5Gf1m/
xUa+2iPLC2nANziVXRJr5cR/kWnWGiG//qqgC1EgG8QuI2YSZR+vl14xBJGE2PIs5p7NNNPz975S
YxQyuKy7QSlm+wwkni0OXcIk5QMHA3tgZhGY3E++okahgABVQ1gE0omeb+IKywl5fLfu0VWMdRBJ
h50JwdjQwIJkgZBjYgqt80a9JxJYsQeA/vZx8dPzR19/5PZ8+zgQ/a7ksvR9fCtDVgAcbOBeXw9E
uWh7xNIhv+T/umV34dyLjhD95wSVyBmNof4kGyO59LVj1lHevvABMZji9vCwYES/ftH85FdGHOTe
okfKv5Vw7x8iyy1p/PKyRZBnZ5hs+Mli5JDHjr7x5KZZC/eN0eII4PBO9tgj8TDFitdLEoSlAlbQ
OF45AWat9Cq/GEitgTPS858OgNU/nrIE3eylqEO4NBq4FJfX0zaK5tlT4yjsFiO7kjAkpM8aHQ23
8f8Z9jXilEXI1f1Gi7Mt8PzFIfVXI1v0gvk6jqg+R1Xpn4Bi4lxi6cCC3MJZZYd5Jqb83Yhna66k
XuOYEW9NLT0dgZ2Ubs/GwbK4QtBYHYmh29LS14xAwzxzdfA1pUAnq6nVrdlaBF0vwJPg+p8J5x2m
TA1rOrq4R136cPHd/TePEZaMPe9f4igbCnQ5RvEE1BK6HK4iZbeKQ5WudQvm0dg5xdN5g9hbtixf
1Blu0zJdHu/Os6f0OrYg/t2uedpAylMxCx9K3xaF6ut/0kxeqJTpTVC6rum6AjLBxG0O8YqSWdCT
Spx9YqQJ6iFgnEEayPmnQXlZlRSEtf698JBUOCItTQwUEe0N+ofIGsOSdZoYvkaDTDjiCUlYNSli
EMbE3N3i76W4g9pGwVt94Leq+ceEmj3rV9PQcNbtsG+UrmMka91CX449EMATAVuAl6xeWaedemxE
VEolNxaqIjYbTHJxJc5JXipY2Iz7heiYd9w4pi7eeSWMzqhtaSRLlWnqQuek1ccVulg0Ff49uVwJ
rSaqfCg0shz1yynA0L3af/FbCTvwBWp7k0iws0SKobDzc3HF3q1E6rRDdhl4yQu9V4bk8tgWAsPE
92Nkk8MMFe37N6dq0J1aQtK6fm+yusNKIsQLJWRUJozvD+qfTLb8wxlAWVJ4fge8k/UggjDURFBs
KRXJ+wZO36vCGQ3Y9PXF1BTd4x8+MlCOBoShvWR4fuOn9vyGdWrgjJhUP61d0aFY6aYXgTLOHryu
rHo6EY0B6Gq1z7OrTUzEprvGDWTwPwtW02DMDShvz7KQLIohfgNW/hUxEA6ZpVZtyqpi6e9VpGBB
rrvd2u2+rrI/fIB6lm6dN57oWDFKczMJV+12ZPOeVLSCJiaer83w39h2qCAZ+CDzXpPVLqyy5SJU
t7DANhBU6W/FhyLJJfo12Pe42ThtHNeIOmJYOIl3XYxKYudbETvAowonSbtDU1aRQCCbjl8JyGpS
nkmkPG6D9BlslNEkfFijG/iGBTk1wFA0O663F/f63Oi+9eUpFmR/EW3v4Yck0LdtHxfYOxUBCmaW
9K01IxB1JLa03h9RX4u/lg2otqoHnTNENIaRLeM3m2mcL6JSQEv7bz7jZFtV315nM5eXPtpPJjzw
+nM4yYlGxFH4SE4aBPos3IH8bGXw7DJBLu1WEDOeQpIAMZgA3NCWpRmMrp7hzk95pocGzp0+JLd2
RFHMjXvWS7DTHW7l8Lc/3WJDXL3ApEsArDYRIZ9seSPHtJzvMeksj28mKIm+w+//qDDVAR3hVO8t
VqDXYwAEkRO0vf3nxqcqGHSFmf2HBm4aXmo9prDZRysNL0SdH0Xh6IU+2Fuq213dexChsAkI+G5+
PLHk3dToTLPRPi5g6fC+sz1/bOB1+UXzgCejBqHINwXXa5B+hgsqsyLjDxnLrHHQLZlKMEIOb1x/
iuMGZD3Ol4FxBNfn5YohPYVpKsLHVOfSzc3ApD4FR92xcLOZTJ7PuMiT1Ej61IOGTyYyLTKnIoRU
tt/VetukJktll0GbzdTFzAZ3N2+E7Cpi0IL4G4tAPhAoZoVjeUQgA44nlxHke+KnQL7iNqQqYV/0
PQ3AV1ihktosaaldlK2bLFPN8MxxB0g2ux8s7NHKzzxXiTJmbMgXx4a9SZtphezjobTmDz+VqaDF
bLIxOBQbXo4iMIj9Ma6hjdOKjgbLA418+Kt09b/BoTeejrAwvzr12CbwzDp436mGTHEJmjZWBn/d
9QOKzHFmGh+/aqRXglTq9SUQ3Yb7vrEFvWqQ2cRzktEBYcqZy1yAIS7m7LcT8NOPo/51OCzhFQon
7F3BUh/ezklWha/w4RmZE5BwLHS6RX1chlNcKkUGp8O9rK9CWsHqdJGIGk3J8ovpMHviyAtpgURA
YoCsiZgq980Un0YkSmCf9CN0O2GvK+gpPZZlPuUmlB+twvQYLGyEstGcjakM48Yyea4ltkn43vMa
v3HRvlk/lqZ0o0xHPA7G44q0bVud1ITIRMo/elY2tLyAFOFHtQXRodbZMQCeFoPcwQLobzrOUVKe
PYggHpOSZpZvJ4Fgkx24Ha5JNO5qxBYZ8odclBCYE09T3Sews77vNhjueWf7s83447EN/PHZwAvq
x6sJrw9gLYZR+lXsX54oXKb1aN9cK8pIoStJbJwg4eWxL1+et5vUhK4rf+jtJnbo7a1RMrw+OhIn
l/CoUjSL4E8085kDhTiSbvxqgyjrQGQ0JPGejlvZWnhOdwtntaAwrZCCL92ywzPWbDxc/gfGHjf/
nNZyLVlyY5qB8Zz0WAogCEyZmg3OCsQbWLhAh5gwUEmnFee2ZvtPPfC91dPKRAe1k2fSSRCxVvxU
KSzVIqFtN2gAyffba8VdBXXRSMC9NzBkVUWU3d1rPGuIfYHme+Ruj2ORG2JgU39KdnbD2p4Rf3+i
IDkjljSyVOuyEwsQHhNl3fT3TlCUO9rxq7pxtZy7BLfibTvWjEQhI3fmCTVN/e64TWX11XQKD5xC
X63u/zIe/0vVzEGuD+5wg2/YEErTgzw7wKSq3gHUjYlAy9gcp3xIBtX5s0+0SWQfLY4WmuXaEMlZ
a8wQ+ZHtsg3nHhgNMzf4wqe9uTQ3d5tYrsSjGMnkvgUHNkoBBvaCKpFXMap4TZxOlHVxf5nLO7wS
wMfGSCbRwiF7NRFgXgOQS7RLXBxkZDP0ubd60NnMyzGrrO10CoRVLm7Ah//TydM9aUKzN5qL5eWp
BKiDb/oz7yKjohSSD2NcONPhIxm9DZO9RkmMgzBcCFL2IKJUyuH667LTpmvGQWdHTD/73D3CbBem
/5GmxiGHvvg8nlspqg1XkrkWsKzNjpNw+tOecrLavX2EyxDQUMQAw9/WWj9XK4ryBM8p4jkhRtfR
zwT/h2IjTdYdcbayTalIym4fojUl0ncJ1qumKlDJ2lmAVI7VImkuQNyZsHCW/KOY7mYvBRDTJ1oB
fDqoTtkPi5tk6sqi513lTEEhrZm0OWzw+1PCSPnFPzPIzVrvX8miWfwW6cy4OcqDunOl6x0X6GGf
+D4Fy89RHNxKSbxVBIpGG8NR/ZDUNdYhLrSXU1uAA9dh7CLcZZ4TZKFfzxEWZUbyWlZeKvrAlueh
wdcbRAQyo1Y+v9W4qc/42UgJAyLxIqKmvus58z5y5EDxW7bVnSmZGDlIobHrZeveNEQqiJ2DRz7/
/Y4uXzbgkMYFl/PWeRjDWkQazCBPOkhciY1x9fOGkEM5dhovgJaJBS7n5HsgVf4zNwLqVpJLRyWD
m8UlyubNZb2Ktlku1RaO1kyGDjaKptk7NCbmQOfeDcQ/AzWUptn4cag1j461TUbQsp23pemTH7b1
4dJ8EsFvQsvMUHbK25rumKOQoJfwEQgxY7hJTOPq+uqLyff2LR5SBpMwKFZT4yiXy3fFispu5JMS
W5MB6w3n2fJ8hCGSVKVpz5bWdLlo3rNhDm7lGxXlvgt9mseviA1PhDo8CZO2pvcPyueJR6wxYs9d
71K8ebPVZqt2OurNTYBJEWhvfQOMETNngn5JWMM9YX3OTU5L0s1kWrrd/uQ6rXvzRDIoo+cfF4EA
s4cDTXdyPfKxkM4mBjcWanb3Qyzzi9NH7vFH0UOfIgA/KwyZWnG4xTMB6S8TlSJOOmrVafPNiEDI
ygW0e6M07VQY7ocp39BVHyDzJ7S6pJ2tlRLHB0Pyepe04fMVziZFyinPjmfSDN5kOQW+O12B8Db2
Z44RmtzakDeQDuqJPi3xHAwuzDFWV4Dyl2gf9C2ASFfbp04M7A2VAZ+cq2LEODfFxRGqnIcWZVET
7Yxz3LiegxGSF1r25nRrXZB5bjZCyMk1qM/3XCpODWYtj8m/LPFzomK97D86PhYheTfsz3kKtpTq
jN6vNcSfsSOZefMrABHnfnVTqZF5MMxHLd0mfSA8u1N4tOEMyZGVNp6E89sBlr9z8K5sEk/pEwlG
lTCn7td35CdqiH49ByfMKq2czMWbWDl5DugB5lxiUtpjVmAuN3l/HIKWej140XAWJ0U0DnXqLfH2
mh1fDg1J6Yld+HWufhT0gk8zh/k7NaH7/9vQCU0cfWxVPwwpAJkq1VyQVRiic07laNOAlDgNuaVW
6JA3ViXbwuydIyMj9eAxbt0q31S2b/XelM/WznnM1XSjB+XtozqChEm/0X+UM+a4ioYrUE5ELcre
rutI7BuYFQWVIhOko6m7pTqeaWPKfAydKU2Kjj80/GaVlLUKBR63inaT6h/8aiGq+XVr9eG4voXz
S7CuGWRnpDw8qqstEpR79TX5QhgbVJs60Dz0I5Z5A2P2JnDHyQ+6iW+RXGSVvQKzJT8KHmFmNkc7
zHCTW5XypTGAA0UDNysEPxZzecCX+VH5pecyGcQHoffNM6yVrK32Ri7C+nSwhckt6BDjvPPJMn/L
oJ566lmSMfRl5MPi0OtGDN8s5Y7QEOBvw6m3kJ+WDL0Vm1qgOdThwVcXUx/v+EDODMumJ7iGbAVb
yh43iOTS4PhO6Rvk8YDHy+TB6zfpCvNdiMBhpjuTJhWHZ2KkgkyoRuvJUU0ArNhGW2qx5mqWDMlt
qieaf4D4Q/GcW8y/Lzs/tc/07CGB+tEju4NY25WSBPvpmzzuwRdsHunCuciW25UROsVKOOq8zJ0z
vCtYDlRnR8ccqaQ1hy7YOvJLOi1rR0Hv8IK4ndxaJM3AAhAOGrYxWqK1duoJsiYWaDqz+EUyxIOm
kJEkQEj7x7hbfVOOE9loE143y6Y2NacqNkvXWRQd2KhY+RR8AtrDI9j/9LyFyNIWTmZHmgF6CrOE
nqptKH2yU73ZOt3zgMiE8hfYEFKbfSCiaNZIyp+5CG4kUg2VfjkkCldVKDLgj4paxIE7dGVImohJ
cVwFf2Vg6bYjc8SADgZzScDVSSGbiC8Aa7ml9fD/oRXa3fDRuevCCdpkAFixcI7AxdI9lbJ1NFrL
WPSoTuXu4E1GQ20qvSZSSN1VopmIcTDBE9vaIaV0D0dW6eF8KTKB+INUWtiJdnRWGATC/BvqzB1l
qtKV7/ggOpj/5zDhHZUS/Nc6+PoINetfTm+CWn1xdQlIr6/pm6obDWfLNx8JXrv2Y2nX91wWnL1q
C31C5wvXUpqKIogBGFAQXqOlyORrI8hvwSdrF3GwfkQHtrsgRpxmu+9h5gsWfgvupI84a93KM7P0
fCa8kcQ0irlwprX5bbHkQ95CllTcQdb7FN70UNhGfD8KMXklpZfClFRcuOn9QDWA7KlV2ADfGMfh
e3kby80aSG/jcsEWeVUvlnn2OidOs7L6ugzdQlT+h4qfc/+RkpP4TYgN/j98yRT8IKXjqODFFERS
bZNRh+2dZavda3Hc3RpjGUwXwCRCXuTuqt93tRsUYfzTpCQdSBWqsJ0q5ROKEpTRiMclIzrLKfsM
EfYTof9obfgdq1x57JtmUNgt0fT3s5j86OM1PWAGHEQkJOSYIe6nCcZkXhM4/onSEVAoQi8e0HPH
gQxuwgkpfUbQ1+g26kRURazXhupoDUlQJkO+9gEw+T2rm6344givc4q1TybrFXyT0L+PV9CIVAiN
mxmgKS5ezDbnL4q0DTnTSV2MOAP8NmXxUU1YjtQXBxvqCLqtMKPbgwuiPdAdGFxxTY2o8tYpgW4u
CDh8wpZY7ld0EGdb1dwzCMhUKDMVb+61gfFpK4AUvZVU5nnfUaJqZg2O/f703WL3+xR2HRRZzHrO
2TWehJh5aJFyIjLFna6ygOHu0l7ASQy4Y4AB2xcA7dNrPlcwp8YXmfTGsx/AvF4roygdiZdFk22F
WfMEnJBJxdSMOBBX3PR0M0sPPtjRA+2aiKK59BTi4SqGsf8B07XHMi+tAAI2K64YB6nUv7tYOJM9
TLkyjYPfXU96+1ldB/sp2rjDdCpMaCelpS8KNVwocp2gphEyvINDyuJ8Hbxpb861rfBTtTufUnC/
n2d/HovtoWdyDltrwWLIhYJY5mv/TgsQOlelUDVecT2TkqCNwubq3fKrCNtKGr/r0rwtCPusOsvW
T7U72FQbsl5HPLxR7zmseheHQHTsNk8kNBkZyzaLWnbhLFU8eIImvtadCDrxdo5yMZm5m/6OSgA2
qOtx+wF1mOABmPVd5bgYH3sxVFaLHnxfTSN8/wqHKGR/bSp3Cc2z6wasn2DF1Tsg8xjOXURoBOOw
Y5XI4/HfGYm4fJhY2hL4kEXbllIcUQSjFPtOMEgOPFn/GeoYlRFaplQA5M1uSVn8ZeOqBfsvKZ/1
sQyvw8DY6Togm0PUeNuxb7ZjHQ55d7SelXOHOHBfOF3H2K2OqBwMVjvvNF9VSmVzClZ1+ElGH1Go
8EXr8s2VK/MtAsNsfTqjJxR/wT2KkqddLWhUSpIDCnRHAKXC//KGwR2GCdWRAuqgxqoFz65eyeeg
nSvVPbuplIv1V+LVdJc6msQZ1QK3JotSCuhA1KiIcsoSGNOEUb+Wdqlo8ws7GKPHlr1jkeLhurhR
F8MYj97cTPaVEZDBOMoxCJv50a8ENjB+IQr3Dl34EjkXTtLXWUxAvu+MFifUI094Kx2V5WkBp16S
22yPDYJOXbHUEouO0+S7BcnmaM+0CJ265j3hTq6bHnZMhuqOcWppu7frmRYEBnwLc4spWsgRjuji
gkkV8MuV7QtINi31mQV6O43CP+OHd/LeUNMUe0Qix8qz4Y0yjgcxuTIfogLpmZxEVZUwniB46cyM
Czhvof2HmGCV5jLebrGrqHLbrdKBGQddtm0VEmG4Q09EbZFAOc36+k/7VpT5qa1Qg5F+3Wc2BMR9
cuKlBAa/QpNghK21ZzG+Vs75Na4mALfchendttpR1omrbrU62jX9fCq8jYRDyJ0EaRWtVZhsR8Ju
FiYTDIGaEClvUX/uAnfWAVCHTdXSL0DdcRm9j0VGMYuYkBWdWKNyACo/THFiirpXLpP5fWs4jDOc
sQ4SfCyqYdKEDFZkjLlwuNgGxkgO+j9nqh2xMvBFxnlcOoNPzuR9qEG/aXxNs36UpRbD2mrxAb+c
PzmaBB6cwO9CgAmH52oLOLb2Jhf9V2zYLOOXSu5hCpSuCwo8aw87S/IXrKUvjSPLhfZvJRpVn4/T
mj7iL0rkuOVDYaCBLWCGVNHjURab9QR9Ldj60g/2MunD9aqZO/48A6940Kd/ya5SzbjCLJhh3GcG
5tjUif4GsK6L/CRozLhJdLmo/46bJ97j+7/wrpEkgo5OGTCoxR9VFUnZvuMZ/tzANzEmLuBATVxy
eY/o0ctBGwIrBErDj8InVN9lLmLvrj6TslVJz4obSUmWapuG6A83wWDI3yD0zU3e6Hr1/to5+2QS
a8/k6UoeiLfcN5tte23qe1ZLycqrT4k8AYc6p593Sg/a36uKwluwQAeew1ENkW5Gma38jItjE8x8
mD1Sc6MsVkQCXLzc4Nu84tQ82UDr+i1Pawdx8CfbCzlFpM35g3xGfZM6S+hADELHVyYrdoMhEzwe
U7osqtwuRl2XnOrs30INZ0O201HBvzUq3AvSnCg2iz0ltGD12zriU0fzcA3M6JJ1cAGy7rHHxGwg
MZ3GmB7JRdPrpkXUmC3e0Z8XRFpqKvyFMx+zbbHAF23zupQJyI6OXw8UwNimQyXHDcszp4pLC0XC
66fPK3mez1Y9HLFw6F0+n2Hgn8zpA7JwLbp1BClDdm/lJtEMCngqAgLOMmJwVF0gFT0qAwM4HouQ
EKQZnbj9j3C+fGVrVDglRDwfIhBp9rLY1FYdoT32hB6N/9JgZE5kk0K9Jzo9wxESvJ5u47i7YWoV
7WnXB+iSyN1v5NUqIRpkxJ0Axkk8Eo9iNvj8aPiXgEYpVk5LbLnO0327Q9XU9up0lCaS33jNptWO
1b1mmdy8WbcSbS4O747tJ5bZU0Jgo7iBRBZQ/4TlIMcoFF/AiiFita95IIoym5XkepGYUl/MVzZQ
JAfAteFtXw4EenM2mkqAoqbR55kyXG1GIH2Dc9Ve8X3I36CB7TifB7gghbGmf1BegdQUtJNlcO2U
04DoOxLACgnYSE7wSUOl+6jiQFv/YahJDp7Sc+zf5w8c//6FLfZ5WPcFCjn1uhdJYv7FaiA3/qQt
sq1FiDH9kCtoivfhEitYnmPsyoyRe1gdRF9bm2PLp6Ji5h2feaYd47Ew+XkhGR/NssotzpHq3/MN
xtGPV7erYGIJjCNXz09+SZMQzamIrupipQ0R5BIYNvnFRKKItHIzmCb9hFY9tg3a6LqwuEfiZi/j
NQ6z+aNd+WcCYC3LDvTmZu9ewXGsZadhFT4iegNO6eMzBDBljfI3XCmdWOIZvkR08mrylR0f5qAe
S0hvU89HquMM/T3VUHdLeoJ1BbIeN7hg8yAozU7f2Jn9+aI/aNQk+QpvezzrxsM7z4nk/LDFAH8a
u1eiMdTVKXmQZbB2A3OmhjwLeR2V8EvieyfEPo3rHWZTuFl9tUoW9Ej1/BeMMcK6kNO+RjxlBBcR
4GTEoPE58spQbOmYGHKMMWfb0OsgN0TQpXrx+jh7ehQmSLNVQ+UlUk0vK8cGCm3AjrIcNXMRsMmn
SVv0x3VowoLEfS4EavwWgo9x5PC9rTGwXeGUrjiMlA7wYAtvaSZGXi0/EfbI8gfYvYpX1Rz/5nC9
QfAQFa2jJTLrdJbecxsIQQ1f49Rkjskj/i+OyjLxci3kg4hQ/KFsMF47pl09tAnmdNNrLSnc+6jF
B5pCDX5+IFscv7EGQT/ez6r/33oMu3LOcLPc94hPW9+w9WlDQ0s/8IG9vj95tja4ffiNy7qUzlKS
R9hdeqlJgHYS1QBxCgBTXN0S03XGzvzHlma8ZKcxHqc2aYzrKwN4KhOnKIKNy/PhE6eXZeS+TJUC
SX5ZrnIWmltgxkabFYhj571nY622Ghr8T7mwF4CK/4nzxwuJ9tgysfMjL3xLnVDv4WsnAdndQYt7
jdhJtcCIrjK+HWpogGyPmBopvPvXIZoVctYcIS3jRrp7ZcUgFE2DrgKWlPnNcCFN6EN6UZGJob5i
CwJsCm2SjGLVwmDhQWH4DzrgGJqQcmFHfOcINotyxxjklTvhHmGTTyEq7w7yWcm/1Gi9dCt/jo0O
uU04bRBeSo3y+BPtJtMiYpKTZmWdfv7kB1aI4iswkSPJ5FtHJ7pFusKWzlsUliV5orGzc+hlzuoj
ckyWFCq9YdlIfFUXrYwgb/VHasLGOLOMy51PUJpfjY/ce/Tr/3daHjdvuWs6HKn3DAGxFsunbsy4
IgZludu4AoG3cj4MSQFpHYeJReZ8bPBZjdnUJ62W9n2ENeF4RsRb3+wb7Y4iLsBvCa/uZNbfpzkt
QJ6Zk+WfgC4wazpaIL4jAP7VWBgDticY3kaeRHRqls4X3h45Fz119YnJtylznhV4XUOAdTC2rXa5
hNYxKYclSkzw3e2bFnrThBMcdi4mRZaPvwkKTS2G5VfuzAvztSOC6vSmq4yOnFLV47KkGVeagohC
ucsLL2oIrCBklOJlZJIvZXR77vel3JBJYz7YybWZaN7g1Py3P2BhiGhSDQoZVwGsGVpq/5rKUgRw
Q8UMrL331KAGHUJJ+Gv7LXeM+bqRO7/4Qrcid0i/RDIipBLgHGeJG0SrbM5epS+Wu/8BiAUpyjn9
JQfR4kZ46OfiWk4gL1WY1afcln4AMtITnZuBJ5INKmzkKSaGsCHgmug+K4BSJ1nvkPMzfhdwgg2j
Z0OlVd1o8WtQ6swoeU7s96C0r44iX+xSuzY5o/47Q2dlhhn50hKWLWfEPPCr7PPwfupci1zKeY6G
eH+Tf03RG2XaWoqQ2THJqg1ReWmLMiTihuNyfnGKMSh9Cxc/kfuRgst9VVtcetjCz/qwS8Diu0gD
nKfksAUbEJA4pEg82h4fKDhkGV3Rpg7CqPohDkTnBABaxnMvJwQm4qhVbWe+SStx922+UFYYd9PD
RxpBm7K+E1U4WCja8SVGfizxydhM2eYHL47znl2hQlyGAyU68t1pERdkFhBcRjug8eJOmxkpfGrH
lzvF0z9cOwyDUelOfvl1nTk8+GcvVR/s9r0J4LLdtNSwPrsWp/H3IWeymEk8u0+9Z7nLZr1q4Dwm
MXnXSVXAALXbRNk5IKi6UPYhhCi4NE3qD+Zga4NrxLFRvkAxQYQwPHwu0J048mmKaee+uGcvKZEo
uop9A9C2VslrdaSEG02qv2+7aIgFjzZd/fVxeecbWMM4dK/uk5vPNViSj98Ahrjk1XsgqSER0t0Z
cIxzkSTYWyGfZwuI+jkcFeQTf7MmOmGjGeZyggN5kWlHbhuja5MTIrYJ1OWvXPI+/WmgFHyoKJEx
psIuwCc/2EjXrmlS+OIGrYfFljdsyDMJoGXqF7xdnpr3du0GYeD7OwNdscKewcRTwDB7/tihoDvS
AiOAkRvJL9Z6a9hRPd75zKk8Qj40TLxK9r+FkHGIRFjcxGkIcZ7H5c+2LQp2uamLL3R8M59qdtso
9iG7/8G038T12ZmWCzGsgVrd0CfT5JtaAnEQGkXscC1anMHRQ12bDOZYyOdj594/ggyVhkfYaPwK
gPBVxokaJitX+jyexh8+oi+DwP/9pOsz2ZccWwLB/0ZgkcQdDY6nwszbe4e0mtx5rFYq/upNZ1al
3UmaKSq3Zc0xniIrsdOj289bLKn1IZTFiPod4la2KRLu6kqULiS9s07u7lZSlE8jIuu1FpaWODDw
3Rl2UrABkrWK0Ioq20wIZbP8gjPpjYUMlMrP5jBXTJWtkNbrOzcdOBs8cp8yYRL13kHdK4mWyylg
gLGrKDB4spDFesBqm0Ulpbvs/xt9ykWHUDf1mZPfyCXRGd1fxQ3f3yy5YuLV4Gane6FFTQ/rClmV
R5g+xmulipwneiT2LlCzIk6c7YxxJ9PXZC44F6RWJ/cfdIDhNIL9WFYUhj1RbXwIdBMOmOpGLHi9
I67APLgNmTrW7mJHDcAo2oF3bNdMi0Q3pIGpUI6D8clwPxO+/69HSlD+DkiO2nPLoPcP+J+kkCgm
SbpBFvFe0Fj8NUrGpLPW94HiR81t+fKkEh87ZXuICRZ8nR5OecmUdrBdasGdjM8ySTgVy1zjBhJJ
zE7rw116r78fWU8ukTIGaWSrxanxdHzmn1RcA1zgaUI82WIVYvlkb/pJWVo80YkRcOL6tCYCIf/r
Rtt6qTwJQgo+0e6PZkK7ganMNbqKKIJuNHj+AAr5aCl3wmji1gvFX3mk9JJ3Qb11AIas+E2RgZON
HGXyhwTNQE+8aUmNCdP8Uc6gjOYaO9oIp36z0ycBpNCKlFJr4+wvyza4HGazCojyNPhxpGzdwrTY
MGz9mQrvS9EfSlw2kD1QPpVvZFx4ak8v/uNLJikAX+G5DgVqupYE6dOzh0wzuMc03y+/QWAQj3GB
3T3Vkj7qT1y2n13IG47TCsOb3WwbZ8AXeinvZCSb07UPysmxUhvo6ekti6qY3Ym9W3NWUX/eSukO
95iIbPK0sBovkXiUtRju0xhkjzrAvWVFkkW226Bup0pHhnN/tYy3A6tcoIBuKYdWTtDDJfmwlFWx
DtKBeaj0CrBVlmtTsbPg1+fxv4mGyZf+yukbIGqlS5R0r7z/PW5xlJyDklOyWqnoA+jA/Qnn2Uz6
Fd9leBj3/gkH+UsOF/xvYpfEYUZXWDf/pC/GvwDhVPhU1nRHVWqNn36nNYC7Hwdd8p+s+VQXTo+X
Kp2c0nflMn4+RVhQRo1pObPRFCZXfPUck+f/D0ICNFclskjZxIBoTBuJh5pBlw46coV+VU6CBtuB
lyLGeoDUP2ojXrq7WlgeSXQa7fVpEOEInEvjODsP8wDQog9yHfqYNXEYGTpJWAwTkvvR07z4ODJR
ozaQmzW8+CQT84Z5Oc63QUGNWIirwEB3JVUpkfut1rYjTbCxnbHF9n5BTCzflqCnB3C8kCDZrIBS
Igdbcq2jucnu9k5I/mmNfD8LUp+DezD81acj0EfPZ6os9QY4yxEz5lWv63G2y7CWD7yIthPrtyvl
d8uvtrnaUZifQTawk+q2TOrniLrm1TR75/5lu+AC3N0LQ5lQTNQwvglRlF1JOzDpY6Bt5+MKxNyf
hP2haGgZVqCZAqqkkD0PEqIbs4VhCyPm3oyJRZtTBn2/xObDbALcT00q+bcpKTgiSK800A46lh0S
fObuErTD/9ua+Sep7Kdt/DFFmohd+cb9zSxZFobX31J8wmJkpNJjsKw1VG6tfLOoPDj68a0Y5Szk
lXWMCpLmOv9Qppp0btiIolHhGcn8lr8suYK/54AIjydnT56RU8CkmVevZlP+5VdmgwzD88XnKlkd
hXvjZ1aTBskq0rJqXX4UaT9Ne6I6jNP7VL/2zcuMFqaO8tCNCjGEFTmJ7IfnMbnWKFI3rnLCsmZG
qlsLikyOEJIW/VykyFczJd+VwWQFvnaPAT+b6ztd7kakarlmjnjVvlcqJWLKT3nVOTpLxy/HdXdb
S9kI0GpOzo8EVSJfIRNo3PsoCUN9vrCNhpDHaGJm7twlazulN6mfdt1yaahtj/RhAUhSvt3MIO7x
Z/OMXe9zat3XOy7A47da4cVBZWgfJWKT3z8xQP4RMNB1r4cri5g0AJXk1v7dgqTtKPIA+wHFrd9h
LiU5D91P7JnxjtNwFgX8xBSwYzOujhYO6zRLBRCdxtE2/OeaSqGwHecXO1lPU6DhoSrfs5RKResb
uc7Rnmt8/mpBvatyKg2883THLwy1BGJcFRhtJpalYSKpIFapNcDEorZggr8TiQLdccf7975OT2C/
xpWQBMGX3V3tMenEdPhSvThfgNfmQNCSmyJu+tiMGlC5B2N6/q5OtUs6D1QsiDX2j5bGqFzV7Udf
NW02WKB4eonCgZQIo+6sqjEcV8czdeYZ/s+4NeX+OFyZlWuUgkdItpVejjRgEoLdc+ekjlGjBYS7
25GOA+P46PQeIztjhKotmSBo+Yb/zHiJFBxENWI9+CaU47s8f6ARqrUKR82trSt22jdIeaZesgbC
xmcVQ2lvjyXFWEjp9LWCqAKfOyK764vBFEQdYPB36JaL2ifPKrV/2AYj6tjViokJLWRe1qn65zFi
rejY6wU2HNy+/AqXTDMZWX+gms5jHMV7qyrdhjN9NzunYEVEHxG7673W14Vln4LBdgEIOZVet+yC
4oLJWeofwpGsNhRPILK5ZJ/rHPBUgYg44YN/MFF6Mk2FlYMc1CzdUUAiJu69CF8RXfXat97hEV7l
lMrc3+WgH/+VwHG8qpno+mmB2QAi5L3jr2KRtJx8wx2huVcAQ1It+YsegqTSW5JOY+inYQsahmxl
UWv5LfEWDDiIr6lmG+1JbxNNo9pKx8fB17VQWPAn2l7c/152wFgukKA4B0cr3QC/hScMT/pM/lEh
qGKIF9j4Bn7JkBofJpPsVjq6yCVKo3esL/G6tTRq6D8eGIgNbJHK4gkeXT2fDhO/VnLoay6DP67D
E6btUxesxb8ttBjaga8gLt9Rc+0qFI7VRsCNj/LjNdGiwF9eiSKyIeoNyCeN1+xL1N+LDBWVTYSE
QR3Ewu9msbY2nY1E7K8vRPtJ7G4Dm4qgC9U1L/C4dCPkvykH++ttG+y1vCjbdGlbVjaG7yTAiPUw
cldiTmUYZYRJYztMnvF+OvE5YFwIsaWqMqENVyr8d6Yx+IGKs9nOK6BxjcgJqBioBGcxT5oBKOnz
JrtDyjeix/mm5UQ4rHppi9XddeqNhWqtR+adqpnp8KRHkpZfZfsacuyO86mesCKhTK19TKy4pMJg
AoDZ3QL94OCa4RGaFNqIwOcGIO+J+Xze8xUebGhTAWlxave+Wmrdh80BidGosyFfyXf1aI+W1Vnm
6X9A/HYp2yeflsqBqTzLp6wGWQ+rn61WIIVdkLp9C7bP1yZkMh9V8+3bJgg/oCOLfw4MvpN4lJqV
p6yWZqxMnEG9OCkRiX+CMjrhDQx36he2SgBabBVWbcmhHR21TTCO+R80pSA0eDuYH+/ZL5vZjQ12
Ai18/BfjrzTuKlwGvMk8e/UNotF7PQ3X8nBGNvHZ4fpG8L7i9Jmo0IGEQEDXoBdyRsU6K3eo7Qg3
ZP4PvwURwAUkebIA4gy4z0ZUL6D/rUPtBvx70674LaW3KckUIyLvN4eMlWEvHZxT4HOISu5PN7dW
Q+9Jh/6csCNh6+HUtamdhqIb8K7qc8+0ykE4wL9dAlrUp+SDWgtEbwxMn9PaHo23L60U70quEhvS
kMM7Gzho7q0khNhCEKL7CPGbfhJ+110vSbuTjCpE2VPVyq3ujHw/F/CmS2go5YrMTTN2snuxWsa7
bTD3l5AGsYDRElHWguMJRGc914S1SMRwHuKlBFdk/bXuAFhfPcS62Obh42o74ttyxthkEK+glSc/
Y3wIJbmrltnzjqd7e8UmLtAGoyzeKVWSsbP9C20UhNBMtYJgiIodUDzgs3tC5inAQs+1LO4kZQ+L
e0cD0+2LwjCJMr/+hxG3d3hKltwnNgvfdI5YcdnSEBfnVLAmLaIsXISmP6nLFs/6x5BfQ9oZqgJo
Ro5Xbkrz40U7vfHfWP5SnhqRmR6kD0gS2axZ0V/yce49ZzwBSgmeOWbnuXoli+CTwSZItq1R2jWU
aWv26shEZ7lISqbn54qxUC6DqAhmbr3p5l/9phpiF9X6ybBd9STKWbnfbNPy/iV9YAkFoPbP+Ylr
EkA4fSYuI7Nlfqo0PN+swsWNRqj0zMmrXW20OcQIG9aOwBNRocKIZ3fQpaHjBT4=
`protect end_protected
