-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Cb8FqSE94IiM9Wc7bWLLUFtjlwc0bZZUx1fKbDSve2sUkp0swYYPaAPQclvPu0qGJ2OMThTwbX/8
ZA3h63LX/zm7kmrvww9EU1hAEncMg/jvK+zklz+AWMnxqPmFrKjUL2i4GE9QdH6IcsRIaOlsMDhz
1f4xhx6E+GL7taHPNYL3blhjg91rYJbZ5m5H1ehc5dR4PkcIdTYyT8QoYZLB4mk7yBf4BT65UNdt
LZ1D/JRTGBeI+2bPIhwsa/xSu5Gm9z8Iu+zYd+UMY1CIHz/U3AXlAGlJOOBFr+gQYWgzhztrok5G
JTr/uJHZAIUHxPqI6zCrKHNNjgLzdIBM9mwqCA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23248)
`protect data_block
I2yNeSVGCcqB2QC9IJCQQnQU+1EfhwORRsXw83o68IiVteg1NOJ+/1sWQ7JQ924Kk6FFvbRIw1AN
RUsDhIopou/43nDI5mEbmRhIJtfzHGkvyvV8jAF5hu9hOlulRLxsuvJa892HZ5ZSzGDsnRyla391
Z4XBpkqQMbauEN06Cr1qO6McJKm8teYaTm95Px/3d9kIg4iadaiRKzoiBDObGQ4g1NIhnQyyXuJv
GgJMI6CQPJIZgTX4YuSOrebiDpaSg46roJ7bMcVJxJZGE4KqYm4Q3v5hzHcFvLNlOZXIWXvGJA/Z
+O6XZwXn0uY9/8S/0zsW8GMTjI3GIy4RegZl3S2uwkro81VM4D/hKEzMNXG3uc/vPV2yuZjfTIPR
UCuawqYZrHBUGvSl7BuXoyJaHscEbofwzZzprAwI7gup3VAAJUFSYQbdOGh1B7gNAwZQlMQV/rL0
h/zM2bptrtVtORG4lfdjCoW1tOWvukVdEbK+Mwm9AfoG48dzwVNYpzwJTQapuH35tSkPCLQrZREP
9rN6W1JV0K+8KZKyXU4Nt2wgXekifuG9tCvolJrKX9HTWlSfBE3SckcCS+lq0yuC8qLfTiYPCjjx
QNM6u0hCcEhfIMrh8urUoN0c7gZI0JINGVPxveqSCCW9/qkDMcxPAST549uP00zLbF2vEvX6aCvu
2f4VN4hv2VCvlRmipFQwUl0JiXxbrEkm11gLVVrankzvAPpgqV2NHNLTk5lTbaYS//uqNVkCUsSh
+corLOh9Re1LZXUziZO9zyKL8lOkA0DKrgVbrlCyqnxml55dHvqxHuIVdsO3lxTo44H9ZyduZOIy
poOYFnV84sFCwk3mUiytiEvkIFtP8IJuKuH+M51qUfYlap/zcg4M3Pvk66Ls0OsZYyD7nIoG9T/T
M7ZQJZOOBW7MW48qkP2ZJEh2fqh5sGrDIBgOE7E2XPIw9sms29PZetgVc118v7zf1SXftNjB1O7S
XdzLDzEU53911WYG5oWaA5pDMGNlbG1wyJVKXL4q4UEJly28tiXFISqZohvHDA0pMajNI/SCCA8E
6akzt1YePMQ/YTH8A96/92qAGkxEPmV4WiNJ+CnxfvWm/WPQWIi1zVAOhQSGR6hb+hPmig263x62
vOavUiyY9FNtL1HyBnukVZRMHJ2+4Xm4VzYxy8aZiCC4fPBddy5JktXpMckB1/fHOKZFPnqiR4ni
4Z+qCM86WjJpMDR02mfB0UkBLb051FtaFb37N8qC/vgOHpXV73vF1MDH5gxpvF7nJM6CQ0pWMg+i
kzg8Pao0T8+S6uyeFsUzANEZVqMnItT3eLvvcdjEv8snib4HEAiV1HSJDQ8rS2AKx86CCHklq3Ky
ZnpBigzdjMOq9K1HKFYAfoSKihiar3ezgyGYEyU0sG9Su18IQB+BXW9llAbygXotBNe76uci+Htr
FnKPXZzq1exLH2qm1JtYqpoccvFaJ74tbN2O30BB3Frqc+/w8yCyTqsEoDBE5m1O3qJ8mtd1JnnO
DcHXWYNSiHqOiVDjMvDFnJV/3gdUWQKgXaZQDn3hRHq3GqH4E7R63b3lXKWgcLBTQ8/AaSYZeKcI
+pPpTz5WKJTxOQA0za9xZ/V9QRqSTzwyB3tvwC3h51r6KB7kXjCkvXuNp3VDizcfB0sAzgepjuvJ
+lBmq75ogu/SQw+GfTRIQIQrCYjhEtr7dKyGFJpogKGyA2KN1aeRQiJpXOHNUiOec20xn4AwAiR7
5DZS1+bA/lnTFwDMJAF1vGH4uG4wy5DDW7upHYYfPW47hw9RCVRdUtJ8I1NW7tUkw3RWzJSgI8wG
a8Oc6p9oheJg65q33/FuoLz/qdgBp4gh1X0tl+RDFa+ynSCYG2me+/N1b4g0J/ViSEx867A1XkDH
MVd95miLNJNCPP4Lol0R4GrYa//i4L1ZHfyBIM6kLXQK8XeOMLq7RMSyaggAz6MnGe3MT6egVO5h
SOXUUDFO2XXrjwoY9MFQ2YS/xEclhCxOdrpX/T9ib7/4cemuESs4Kzxw1ta+r5bpumZWgSqqy/Gk
+MJm2tOb9Vb6+YiBmn/82P+nfdAdvs4RBTRv1Pr/vwfF8hcKZ6Cpwuj3kV7IoDt2aykb1QeboVqB
MmtoiM++bb4Ldqs3FnVaP/gad4IlDv+u/BGbjvuQiASUQj2fXU6cdLOF7bPnbzU8ZNq8XTYhI/HM
AOFa5ZJfe29v2TA/SCDRSWib1oYNM27N1V8Olo+Sy04m7zNvnCb8FbgHdR8BlfFajdQSPSRGPd1G
LbXdxdPZOlciHnyTzB/Fry0lYgoxthW3IWihYjHbEjNCq+dhgbb4o/ZHWcSjmoZrlwGKxdfs/PY5
+p8IV2bYQ0hCfhXnsY45VScOfjkKYh3bACOjXQvFNexxXEqx2mokHI59xHBCCIZIIQnVyyGfnhvW
Pj/njVCt+h2aBuf7x6YCkFzRx7WsbrT3im9LsUvRsxhhLpcyaDBfTYRw83BSt8CeF4V4Vtficfck
CzDViUM1Sr0zshdHXZL8dNcfsm0SsnypubVNP1YSdDU3C2VwVLErpJZAXzYzfXW2vcXOCW25HkRp
Q6tFgwBI2kbp9W60axUoEjzQZHckLQlMJk5ga1DC6kG4vnS+9JKdeSvpVJmOKz65S8IGDU39CxIW
ClNivbvOc8uadjZYiPpKzn9QK8EFb+WOP+w5goUtNUzA0OyMagsbWRylcmt7pmEG/0SMzd4d+pyl
PGLyMZoie6UfQZ+SO8S1n0xIQ89CsveBmQtsz4FRaOQX8vtX8ZG8zZgGWH1zgBvbqgWgOdz/q7H0
MXT5KhCNyC4faVVTBKPJ0Nzo9Xk33ySvicH8NGEUo/MUUESDCpq16qvSbuxsMIbZn1n/VuVw9zRp
qEJ6iQNCXeSx+dAsF2CB0QuJSAxqJgVEouVf1+VzfA5boRVUIa4Em/NLEVPccFIN8JGYE0owx27T
Fj/V3idMkoRaXQUzyrGcdOIdZOAyVg/trwGcte7eto10IJWy1TemndfMAQ62zIV7v77ZK3jCHr+4
Zzxh0uzVOhhwpT9oEh86WnErTvvYUm5T5aPLknnCZE40jgLwJuMI42ShOPHSL1XvnNS4QiNilmUC
zsz6owEHfX7Tn0CIld6BeRh0EfUGY1WJnuTro78EdBy/QcVC1lnJlCC5arG8JroTurdDXATEI1O3
xwsAkwUbIs2ifPk6kv0PQmUvus0bXq2KCnwoum+5SuIHtKrvR6tta/fCprIN1CEFpMWd05LHcDmH
Ylo09PT5keX7et5AYWGretmnXFNAAG8pNEUGA3fBWS/3WIX0XvLMWlmsJQP2Y7G+rN/Lna8hhM38
TJuUUuC1fMFnoFKIbXU7RGvaj1pWPSnekhc24cztgmK432TJ3BcAtFqXQXqHAxVWThRBi6zoBHGp
IplJEzibTLyKcPo/MQGxSMkhk86Ikrb4kLApmSboj2M0JH/TZqqGPeraa5q/OHahs5hNrp6b3kPr
AiJ9PyHBbb9NPiSVyuOw6mNfdNPNCL/kjmx86o0rk7CczzW4w5Fegrx8z0957vMkZ6eDEifA6llV
Bpn4U/zxu6afbjq6hXPkZsW3VJFRHJIt1QXoOYamCUVv3EWwCk0tXcXW6QT+YY0lIF3GuknDLyPB
yaUKTJJKjryQO67Hla3PdidD9UaFOBf+Os4UlNMAfpY/VWjZuHWHIYmBKdL9Fg1SCEHFckW7IwZf
IEkffpDJ0pjrFI4TWGv/0C0tLsG2WunbHbvbDX7pPjb7Snar5G8AWNZu/4gI81Y0JUIdQgNegNp+
JDZwQR7hykd9EQ2obnD9FTGnhPMO8FLinZgu+2I7MkuLWbiu3uiTV0FIgVLzmwY1DSow6JnJxqAC
pzNXFEvilVXVnuH6ftncH/W7Dlkgy05BRGy+HC7ifC+ucu5Rldn7tA2wx9dSG2pi7xYY6IskAKTq
BiWMV4IUkiwzjTak+pHqk9fSueRyJepPeWH5WJ/Ynrf7Q1NatGqWd8VFebL+00GjGZGbUCEFn/+f
c49uF6SmZEvYVW7iBCXRCJg5qqUrsWTxAMiZy4dWWuYF+usIZbtcVqpgQK5ihdVqq3lsUSp4UAwM
cxjg4eWpy4RmRLvXvhmPOz4EmJstF0TAZ/QCGvH5fGgy8gUVTJstgQdjHEWlsoBassUqbtFGH9SQ
M8n6qtZ364495axIMaiQwl48r0z9VyztXS9lDgsYPstRjLizQVgDfwwGaXtBVyU13a2+fF9e2mmZ
Hi94z2WN/5bxj4usDyqGTi+2N3VHe2GAkQgzB/KH7J/Z+DHqPVL+aRT25tTWTs0xPwAlLZhVJQKC
h8nvS/NQKm/R7oM3juc4IV3S1dEvMtXSES0yl1aakM2xy8/IFddFyNGEnMxd6UN9SKHztoE67t7p
vANuCmNyxqQde8wesFDRSI0QuyINjqoeDsgQpBfEW84VMt7l2msh70LEYG91LVInVtBkGvJ5XD3R
ahbBS/kyO0rNYbcUc8hMhudM4BdxY2WvcqU3w9K3tjakrfG/NKIoow/mNTa2sMJahVyhPHuYq5jQ
0gquj43zBDvVwOHD3RJzp4UisdmDrqyE8MzwmOsBnalzztPd4oiWW9VAZ6tJoMfnOmwr4wc5AZMb
YRHkc8WmeFtB6/fuUDvif5B1M0FTFZBshhMU65Wo7O3X5yktcoM9B+3QOclj1k54nxlc9oNSO/5S
aIIADjdRPX0hIH5NAdTHMbck27l+ocv926r5ZbPu66Gh0eJtt3/CUKmhqSMsCli/RUiXIqbwMIgl
OiRSKMvQ9T0XaihfC5itx6TNvq2aMWxDe5bpf5oXQxfCUA+LbzJ5W5dLT1t6e84nuLt6/LXMWRMY
Ii/5zrofxNAt3W01OxWHYgRy8gLymdrnKwVlYfvwuKle5pHjXjxDI8gWmn6PqomPYdXYrRaWe3qG
2iKU7FDdmfuPDDfi1wWN1mNpVkgMna1KtWLBV1nZ5WP7p1xU7+uF/ZlIBncX0zyeq2L00iowm41Q
nTDhBxO2bhZ7yHzM8qDY/f1G6zDZJXYle3UuCazkNR7yePDzyQkwPxakTFcIBCf6osPm//rk4dBd
ikKQTwe+bjsqOHo4XnQQqLQT76hG8EftnV/YEddQxTh/iN/WdGkcWxMKwoTtszP716dVD7XzmiuA
uab6H1FbE6G7v/dpYOokJXxLFHL5fMW07yUxyZ1vPdcUfIFgzVFEGIbiI27LWThaUgofmGL7Octg
I/69GGTwLKtXYCpyNmi52kh9p4NJznbDIOIoZJApQVHSg1cihvF6G+28Hg1PDlRTLoyXKA8Qx9Gt
ZIKsWJUzN65ufYedEe+o5YjwrSDY1yo7b3MlJqbIa3vLp9oyB70u8XnXrvdiuYaulNRPyBm/c3EO
e5zs/F5QCygDiPk0wQ5dL8j9LS8tWCaVLaAjEJdo5JLn4zSYS3XfdtlHPRTz5l0p17JhPW8kOd88
dWAvEyESerpdChfsb+dHjqH2iNBDTcjW2qaVjwn/PUmyqYWc3QExpDLjWvOPwElIH8j+Sz2ncI/X
6e1J860+kyVnSV/+eiu0VVI15LSZe6GwTg9n5Xckis/445qA8BMEST+IiEdi52hRn8LgxLUwGI1v
btH0FnRFnWBShqLvRoMQg1jTpwN06feWrwewucCzwnA0yH2wXqivsooaBedgQAX9lU3ENiTN/T+Z
RkMnkLL8anUzyHVNbIw6a79+MU1m7zdmHf3t4l79s5nGmFhx7CzDYWwNS2eXvptdmqt9MDLSUe1E
bk/BKGQj6L22bYwusuvgGsg9JFtzU/fBgPjclRZ34VMjBgN2eEew361F5G37/ZR9Miimzm0jKB9O
TV5YmntbAjaA1MBOIkbw7rNjh3vQuuDkuErzYSNNCV2LAFB031NPmIH0l6b/J9oCxLX0IdE5NDJ+
rdx9HzQ03kEZ+A7ohfh3t4uXMTqFYJmnmVIrTvf2/H8s9dsCwbS+Mk/fkiImzPYGL4N41Pnf79Vp
dMA22hxS6333YmNZJcqsvOvTkndWv/y1RwH+CQ9cUAHBvG30p6mY4MLkP7FBU1pUvFTs+TiBLW2E
qRQSkMKq5qbCo1RP7r0I6gdZKeELBUT0aDJy361ZUpyc9uua8J1JcTnm+q2i+jx38qf6oU5C3S35
H+X2sbfNEQEsIODKN8xCWnsbTmcokasDvKKbiflpjiP3++6nrJqu8/xleGIcmJn3Xt2B9ClQpfMw
dmFEGGaw69EOsAvWD/2fZme5QHt/dYZFPTZt4Aakz0hqjcJzLKqWSMVynlFy9L3/Hnjx8jJ4108X
GppaTNfJgyus5Ps0Iv3rAT7IE0fRbOgBi2s3szZ20Ya8UTTZZbub56OJwXQx+xnXSPGoYUwmiYSU
bqJ87gZWSio2QNkrVzy5Afgts/ueTGmjFcN/HO9VinygjF2PvHPbQtEidUXsYgt6SWLlBMoaxZe8
rs0NEeFEQdvoFQf4Xv8Gcu+UiFcGuM4PvV/LQhGuopQvk/hG18KkGT0MKDraBGV5gZWwZQ+OoYiQ
YWEkNsKEy4B4v6HlSJUwKsg2ZFBGXwaKoFvTXUEf968AItlQAa+3oIcw3PVcgSg8dWD8VkxXMAuh
Wsxmesge8kVI5r8EhibOZ2z33EFdGL106vfw22TWqdry7j5AkcKvvb1TFfkSPdJRTOVx5NPEoT+z
rY9XYf4vVWW7V8J6bw60v40KuqNzU0QIVKk+8njt/jeL6pw8DCiIeWJRepPCJWU4BKnXWZNC+Uf5
7sgFwf4sQeSaVaSG+1aI3rNewN00pUuCNSmmNBhKq6o0km50CRGxWSpoj3S21MZrcuxpOvEXPLA+
nh3swXRp2S7bar3pxezzOHD7aJ5DqkjceT7OZJ+1x7pdjaH+V8zfuPyW5lja2Tx1BXq3UBtsTZ3Z
cVWpxX5pHeiN0P6ihXNpIjjnJ6oh/55TeiR1bQi3b5rOApvfIW1awIuVL8Vpzg+7/ZEFe9+1gB9O
PPA0RAEtmEiibc+JCN167Y5JswqGrmkBNsSdnyHqJnHo8+IO0+XxTZNYUK5ZMR+V3bw6GepgZDYk
ri8aR+Ycs888UoKJZL5MMvTD3Qbsoy0dltTtyCEM136J/G2rSnaG/FjciMD8+D14pbYg0IgK5anh
vt8Jef4qXWO2rpitUhEtby0oHdAXz5fhvn6OgGpXGfhihpgBVUDZeFCbS+nktSvklcNNE84A8VFX
pfOspPjsr0EN4sWhWnzVu1/RmVQzwtmuvI0PCAim25nf4X8dONA4zzaPEZKHsvAw+6ejU0ExY7fy
TxMjkofF9rzmPQBL3j6OjKjBLFEFTS5pVbUiRTBR0IdnnUpE3euwnrvUTV1YgAC7/LF8L+qA+9Lt
h9Mx686g8jbBMAIIrEltE1zSuXeWEV5Ka0vvCcU335lvsV+H7uov7ZukFMoJTUUMOwn8vR0WCVAH
ewoXXZTQRUPlWeM+VHzdz51/d4+yHksInCjoupVZjmCGcZeGKYXBZ19HSnUbUS7gDixUi7jpKliI
ItKfZgo83R1OJVzqo6+mBu+ZFi7P+O437vI08jG1MrLIZFQ54PhlbH7SCuYnTVLC8F914+qOdlmo
9nAvmbuCcyJXqRkP/lcopPlzNN6Ga/kUfQM9NgCzsYdbd8NdR3JwRoxytf6jhMde/AT+vnmeU0E1
n6u2NHFWkrZOJ5G+fvCD1/bNLTeO/3NKoIp3qy04JCJmN/gFR538YKsl49fatRWfUx3BQChbZtGb
SlFgAqL56kyZ+ijU4OLrJ9gY2kk/2HHIuNgr+6ONc1/MejAb/aYRdPxcbHVPJ1beGgbEmCfGtut6
UJ7mYXN8/DVlEzTnzfl+ZEXtHNcgg6iouhfQJolCOsEGDrdZ6wCmvDywwCciYekrmjwDLLpNUd94
QUJfX2KGZ1bwfU5U2vDGmlIZwt+tNmILKp1oXo9jIwC9A5SSis2EsmIZj6u3nB9kCwXfk2hRpk1c
RDQinTO7TfYwUv7IyeY0hBJ+WRDmnZLUNsMf7B1KFHT90BiOJKmtAbR72WMmfBC8OIATMLpMtEQL
lD5JzxQVcsac3B63bb/T8b6C4SIoP0zpW+yfAKTkI1J4eEiSWIO1zq0Eo4L3wcQ1HwkT4zSy29kp
3jpM2Fpt55Gw30b33gYoWB8X93hMzFBjz7PVUyftDE3pqdGe4Y/UyOBLHRintHbWZpJ1MlnR5mWn
0gVnyDIPOrR7BRVGKlZCmQldOK9e1c29z4ic4XPzRqNdGT1kq29cTtToUWuW8e9BcLlzp/VXFEWT
k6000kajo6by+e7/ivvKek0zsnvXJ+IBJSCjJhpn6+OwLEbdGDpQa0u7c+jRPU/QemO1bV2Lhnil
rMiMRSr+YCOY6jjyvisSt511lcV/RcNy/obzLImJDcZO9tYtrurtU0jqcmSjVByQsEjZCssgOciL
Dycq8JvMqAcEE5H0WhiHeeh38xo4fDhzvVZF+bSvrcEAb5+f8FKpUmFZ9ri2Gr02HQJKEiS+C0yl
WcfziN5y3ZqYZZxN2vza3RjXZEsAXktIm/QmCVX72uE9YxkixqdVGUP99hJGdYQN8nsV5djoXzAl
YJQ7pGiCq+vtY876nBPlwkvLQNnoQtc/rAEfS7gvka5Qc45j+bNIMePGhz40y2D9DxNgLYuSJ9u3
/v+l55uszUGP2AINkz47RHyd39wOFU9Vy85N1KLzKqrScsoAmpwWJ7xYzgJR25ZGSOQzjAbdfW6A
n6ypiljXCyvq5svo3RuibP9iiXmDFQaivLvO4NMBb8Xx137/jCN9j7iZ7bON8Oj+AI8RD8iek40E
E+XGHhGo4ypmGfGdN2upcKDXAU/VsjxYH496QsQEF0iYIBN9DiodIVcqks+CIOGAI8T9r81CH/lI
pzMM74v3AwYUd2T3/KmzR46opli796RbTgncjdLQsperlj8p9mn3bF90TUoRpzYL61CpW2jB33ca
uIiHM1k45fyY/Z8Qln7qz05BElgW/B+4M/e1o/JP02UAU7yom+CFX44EEgxwez/HTVhpOaK2w/F5
D22AxiWnHJ+LCm55sAr7hvW2ssyYKaFBJmV5jEQSNPAyyyJNpmN2dD5wXyyhJ3fkuOX62a7zkxYV
HONZpNO02fbc9L5ryOAIdyRBaCnv4olM79/YbJKjhdBup/L5vH4XzC5INqwtt+Jgu2uJp2aZ5mIV
ghFDvbhwee1VyFNKHzHWaciHlrxZbRoo4AX8h89tPoYmHYESM/xCrV9HHqFQr/r32MJi4HgV1QSo
Va1BVmVvrEQNVxvQXL24YPtlbpPYtjoluO2vVUxnvR2YGe+kcgxD2HHSq/kWrGgL2L4+caqLlMe3
Q8QtH856lfgGij1boV5xW25vT1u2ajzkKZHVYhuEKFaeMva2gb0Nf3DbkVUftxUIXHxwlvNPNvAP
ocg/7rhzmXFQqwRSCqXMKeuzkNbIoIpnCfVMtu3TCs3FpLVsbtPOEA5ULkRMjR1WpWDFzxttBVwq
g5zTE00ev7Sv2xWCdcbcuV7C/sZiHMu4jnRiawwn1kORyWwyb7R2c14BXiBZPFsgvm/hB0EjcXCY
Z3JxP+CsMwgBE7YIg76JkIhhZIcgYyRNmKRaa4o/sRDXtDEK6KqXif39Y/HukNKJ81sehc+AXQVl
MzfbNSWr+oWszT1R6cE3ez0HvQYOxJ+3yLYtU//4nAGHLMoAOEPuNeURoRyR5uY1Z2WgQzB3u4+3
vGlSYQD1K3F1J+qgu+QcAA0085EGi2d8XkS+aXKPoMUCQ1DUFJ9+Pb653TsHvVpHYgQN24DXlhwg
NSvU+a5ofc5VM5XPlPJVOf/P90X8LFkLR0PNK4z/15SPwOGP2Ti23iJP+0uNa9AV1HcqQsCgb+3e
KdVRCZDwxIF6siPQyYzUMG/Q8uqifhSjhIU0IKYqZ1Wgz0x5OFty86B349NcFn1aVtatSmFLa+P7
kzq47wa6KoIEoFerVzp/J+GWFq8YQY7l+MHl9C0hONKPEbqeLBO6GSQdicz67Ffu7/qCbYIqLqA/
zjmPADp7FEUf8E9bivria/sZseNGaIcThlykTEoJC3DeG3D/e/mvhYCf6WqO4Tp8+YLpjnYDjfss
wH2EoKsl+QAiO1IGDESu4diLSjR+wESG8EqRF9jml8MvT3jBAPeqTAq2fiGasEco6mowZtfbTpC9
81tdt7SBXuPJvP53m4SWdAFnAF2tKiWcy3SUgHYReAsh3FjKuapc3dZ9l3N73U5b5d8yOHRMt7c8
o7WzgVkl2BjFIydOMkyDYP9kLnKC2nYE6lchZCmREa8AblPBABl5RQKYsjeMmrkD2W8E1DEMH9Uf
iWTgmeZ9VkpagOFy84H7VQRRxTDiC3zTxani/4lpSnaa1ifqEAI6MtBHH1HuNQ0thhe7dWwltkni
xT2sXZPiKCDIrJZA6K/90I1LclJ3eXAdntvTa/mZKJebA7dqiATlDSfdCOXL5EOUEL7xoNqmQt/B
S4jr4mSIk8xRrTp7kVJIuTqq/DYQAU5j7mbRaBvDKAfdhKmZ6jBRIwwGt1gxAcYDJ16QF93hH3bf
cQEcgVF3EAV0lN4TVyCNtkgR1guEfSFehB3x6xyzxLx0M7htsKyo9NDVItPurTbVMa/MTmvs+DRP
Pp5/5PtPtyFjVIfEalFkySpXqHKGojRYke6UDjHmTaOKo9RU6GGZlA09NnX6GMsIBSZ+n7CSi2DO
V9OIyG7jnhtjuMJCdPgv1rfCFlMXGSEUoBixfyEO+wVJwCf/7iYxWIw+9ky6ufk/+sS79eMZIL4m
hbU0P4pTaW2onKC3iA8eBQtl53fArGdfgrVfB7SlfKlwAnm/2cF9VjIGGqiB46US2/2ZM44dsK7n
bu8jfgwiMYJrxWYfH2pTqJQGdimqKyLuvZLU2Em0nqDTzeBJwbArKjik5ESqCOjkD+8rdTmeh9pQ
Voj/zpdVTqnozgFNCWZeQI+PF4PbsyZOkXLbnlCYq9DcwTCtlfPv9ahY6w+XVGU6HaP0r8EHQflc
+etULeLGYc2xuLPj4T1Kwp7gtPFwRkuj9fp+nIeMfo9naADKV61mcy3BBrPIzaI52gSsn8aKaRNc
NO8iRX1qeWa3AR/ozjXfH3JG+A02pN8VI0GVvWwHC2s31SP5XIGcFAXXrnSGKQx+Fj9Oa+n4TPGi
WzTiztCaGkA2IBkf2qE1WTaW5vy9yJ9WdUIZhV9LzYx2oxu4mluV8xg087do73pingZtom5lRW5J
yxzvvt8Q7enmFshB+YdRl3Fqgt73VfJ6kaflfCwoRN9bWkSkdWzIb+eXzgQXVszEDlJ0if3kT+0U
4Q3z6u9DZIZ2AiCwYxgXRG39GAvPeWGXQdkCIv9vLsqBWFkFKngEdmx6jXWNQUSoIzKWAr6huHTA
5FIKtjEaCOE1Kh/JwoFNl6ks0HDThKg2mkNIZrzc7qtT8zrPfF8C5dYL3Kroxj9Lb8n0S8MlrSz+
REm1GXAROgxT9aaME36zqbOfeX7W69KlhcoUjYdOCMnU61XQVaQ+uvwhS0BgFO8UJSZcaxjuUxKg
yUuwJsWTIqkokWIf6duVDmfFpos7yrSyJ3KoZncOA11h7LfPTGXPbQGudIVWRDwh8MzRBvlnTje5
UxXFv5hVnUh4dqhQjn1KpZxTfzw4nUHY0M2ir6dkV3EwlZQnyxsEy7MNrY7E/Yhf7FbtySdfumNV
c+3a6kYNUvI6hrNc/sSOgtAO1R/dumeVS/+LdG5rqntrr3iiYWOlAowcNtWTiZfOZh+tf7YGDBBh
gvmfulniFDB/njvondrSnmHpFiYZlGnGd2V47cycm8Jyw8g4V3ntResv4132tn7s0S8VdxMknnnt
mGjxcVuVS8NKGlCfX4d64i8kpdp63Zd6Dx4DMQZ1O8Xjo6BEPMCMnXWazXz6x/db/3m2sofgCsPl
L79vbndohYN/t58r9I42MLahF0Z4Za7gYNIem4tGhZHtV4NcPJLUfuxX0WXZp1bImgMRRyNRBdM1
MsuGn/ACR4mh2kTXx1FzHTC4g2pgf/KdwAqxW5ABMv70nt0GE3qkRNsGHd00LWQs5SvAyNWTilMz
eE7WIxOJjdFc+nWGhjNUq+W0CG6O/e5I2bj2fltn6PNJ2D8L33vavNtyL+LhzY9dhbUrzmAumVsp
0YHMRHLZPU/XXDmkYIIH2e1zVdK+P/8DF6nzvOa1RSp91zs/LvoFGGBlOrAXGGvy/pZwdMhzQ9cX
IVwfCMNYq8stKLUrNnSZlMYDD3m7J0d8V6k4qR/3Z0autdddyUTDishTXkTj3UsCPmWDe+p7+DLh
0+nH2d+vl57i204Jqa4c4ZITRLFcA4wD+vs8yCPWabkzVzrVGRCOKTbIiCLAoW0oHexI+yP7FYyG
HhzHTY2E8p892ip33iLCrUo8p1mnd/m4R9SpK04nMonwvbpdsVQvPeQYvXNqpsakN9Rhvp7AiGDC
uufI3xvYQ2ahGo7CwvCV/BtJutwkS4/dvIQyYyXGDInE7db2BmLLzwAPAxGCD4Q5K44qxglSlbwt
nne/FR9dj3p2m6BNlJ3VaiI/iuELxcDz0A7sgF2DH7Mar41Q8txb+9+XSgwBI/8KeQs/915xT55n
enh69W3EsVEKiST7xnina88M2r5HpQnQxsP9tZWxR6cyi/yT4YIZC8V+3RTOsggHd9i6WiQS+WE2
LYn2gNAv8j0i5GW12Q6QrjV8S7RzuKJakNULCW/otlVUL/D3++Bb8lyOUAuhb8yq1FMRKF/Hebj/
ljCzs9JlBgpeVxe/befgeKTPhZOmYfvbzNSpbwDlu8q9/mWNF+e8u1rkwVD6TGt7GVFxMWQ2gr00
KlNexate7nb7/zdXRCRgfLeR98dDVmetI5z6dpUhDXrXLudg0OT/vTgsnAXriNMegEN663grNsxP
vcFgHgo9dP/iNkVI0KGnf1BK3V44EYa7ww3hR4t5oROLH98nTrpgi6145GDW0s8EJ4nYgxE6xx2r
mcO9pLjNi2o2UZNX/PN3t8x0Fcf4fnarZwOQrOLdVOoKa63Ogwz74ksCeHW7duvKcQcDTg6HxG5i
eFGzAWDzT2n3E8SrO9sfybUSBc5dbHPfxiY1vy65osmrqadL6V4ZfypMjkrtaNFnkw/GasYQ+PNR
QL6t5+CUJJZ1ar4WqHkPwByujXmPsCnYNhIAQQn9SV5RRUvRBq27NFnibmleOQYSRu/Q/Nl9efKy
kFyvneSY2LuU1I21zYG8BucWu6CzyrcyLi+zO8AFg6QsK9SAZu4TXK614XM8WLq+4pprc0xYjVm0
al6Ho+SRmthMSMGHs5lkE1Qd9q9nqTJSc54ZVCZY2CHfX4wLbQkLx/VMor0xPMXRiCSl+FSylLI8
qZaLGESEAxHMrdKiv6gedUJX/cHjzfaHZIM42sB3XIHH+QCaUGNWMU6MgAVKL0HpfPbIgEefXah5
RZ9Rv8wEIqS8HtklaeqSoqgwDq+NwKDVxKKUxg2t3Uk2RGyssIxWiJLdzlybk3BIHq3EiXrIrG1t
/w+te4nJO1nB6+Hfbb7mIA4apx9PTLYlkiQZqHbZJugNOfXt+vybgeb5HwGfp+U6mQwI9YikV3yM
4Gcp4HvFK2j0ZCXOwNXegE6dimHMuQxYX9Qm6KcIQthbk/qASypvbuqbNncbpKeMj9pa0XkNzVP/
36i1dpLEEC18tzAhUEMfMFmxG4od0LvJcEhs1bUwAp5WBssJHUWc7g5UOo87meoRbyiXuTDO31Yw
uVpm196f3BdKttKSY1d5a873vT6O+bWQ8dm4yacifqkBmh4p1IdVfupvyFgDFfh/agLIehDU8glo
n8ESnyhbyDggrbEguHSNKRK206YEbzetgLRBuG4OZUPrbAO8rih93brqjIdABY9wUOJv0wx1IGWZ
oeKJ2K98fWsX+1BywewE/xiSb05uuFt9d7So4lzrTHEkJW5V9aT7ozoCU5lAPEwNT+37bjCbmD8g
K1cgUAiJpyW+HyYvANEyYz06mtpt2tpIi7EPvIPC5OzQRycNg1JjNRhNzp2XI6TCYixgEt1zEhga
BuTdj+j1yGH1hhzaeYmUYU87qcXkojFJHUevDqM86UtD6ojEuAsrq3F/AJCIrRzGVvbrVcsVPMM/
lueO5h3Lxt3s3rtpp2DCzjzDBb9hbl87IRgQcA2u8GXD1HOyes/EW3zlUW3ftUqOML8AToCRwYiT
h8lN0eK98Dl3DuijXyBvdqzO7hkvQC2td3UwwlKj6eB8hq42EcChOC+52p3bf4Sl7ISDOtSdsUo3
waKaOIYWBYO+P1XdgvHPcJNyjD8UeohA2U4AZ6baFOhV9z2gJlqfZAdVYrlJW6OsgKEasgA2qf+S
cDr+4+E4zR4yjH2qugPep10CUx7clL9VHPhiVuS6WU5sblXHuk1MZ7bssQEd+swqUMA4FIhQlva2
XI37gjyLeFztd9C64VRrCqCMFyLgTX8uF70nlNlgZe0Q9h/Fbn7ensDkjtCH96orZ052CJXbVy7D
A3eEbqevjzeV6Gn9DLiFG3Vs9UszpEbv/4HbS2V7mapS30k/dz7gOvA2oPjxLwKRXvxsjTt/rApy
ywemR6RItiytuvH+/U0fLxp21rJ7rfqCQv/kw2suupetD4KEuvSPbGEhtgomzaPlP9Wv2rjPdwEi
DzXB+z4zJXlRNeLaZwFH9JOy2J5zFIe2QokoaNyGo1LD1XUNbsdC1DxMHuLB+UG0zCRmJ8y7eMJR
YqEosXp2gPVNw3jwIWy0ET6ggkUx3U/L7qIGdPzRPxSDWoUVO3Q8PmJRa0AMDaHOrc9QNPqEpM9p
ZiyLPvlwhEPDf3cH+SNOhIdrcTsgeLVmG8v3O+5T7K84TM1S5XNxLfiX380/KtLUHmP3eNbRcnk0
OIWe2OiEQ5iOtArKPXFXiSYpX/0WHgtfDSbwgq/wmkBsuPcJgnk0ZTYu9oJ2VOMT1ouO+bJ3hHew
miRC1MDYKBX5cmoihrq3RNAB+oANqxoKYmuaxNtjLTm2WH71M5/NlJQDo+tpYS/HyuXbfYMMNfXj
/bRDbycAs00Dj0rZDP3vVwK2vIPuasMs2WQrbyV5RpAzYp5Id+5BwuIFJpfo1uol3AHzwl+HEoVf
wi3s0QGZ/MBQuenZwA3e2VvMt9vRqMmhwuW9ikeD0uQyKAci0+U9ZRufK1tg0j9XIGAyfs58+aSx
dZ+VzulFbp2qZC1iHvCqIvZMYf4vP1GtuyvbDMPJYKYwBv0B+nn9gikwujO73BC2PjKf46VslKgz
f+SeiVVEP7Wbp5ZShHE/5dd4u4ZrK5eci/kBvzJ3prYARRfMF2q1bHSygwlFngm0jBbiPV0/8b7b
Ast9QrCc31mgllK66GnGUo4vxYvReYHM9ZXuI7VPOLoWmG2ufspFL49TVFHhjmtmfHGNsXUlxaQp
GbOFZ5dasaUuVs2XZ/U1LatjlWSZzxhJvP4XyKtIqWtZAZ76cYQoGwZofsLcaFvgfbnTVvtqeZ3W
eU6bZ1e4BBEBNtGDfi0OCmmTYAJvDHGfjT7Edg0E4ZF5mNat6/hULD53/ljredmxdGvALoPYuWZi
Khp4Ko32Zqfh8dLE/cEgBiYwFpQSJzKQFLweARWJLgri+Ak4PPMKCwqeS+N/B6xuNl+qyDOVcMWW
yBEZlycy4SnbWYg1kSqOuvROEAxNZcQ5R8/2FSp2L/cU14ZehKcz48W4iyY1okAljA0l6Qr4B+gL
wOL10mQKVXjULhIaLSJGZOk9z3H/1vXgR3QrNw6e6UH4c+HAiHX1JaOmdBhKjKNmc9jXzwSftlyw
hS0yFKQ/YRsYQRBgyLDVmxXG1kk8rtduT9UO7edfDZellXyv0jgS8kclcA0IxcWDaadpvGL5JM8H
tpKZ4wi689uiDdlGNnYqhAQQoASRuxo53h4Vi/zKvYHe3bnRV2rTrJt7VGwHkip7OnrpV/DfzCdL
RU2h34CLlMdm8TRqnSL/V5g8yAxJH9+bINW880ADdZu41Qtv0nsZQCq8wB4XIFFWbiNPCi+EodcO
spFyXxtHTTfddKuhDZt+0BHqukshXLUk3WfVRVjMM1AcemiY6ajrBVQNaRyFfxorwP86t3KZPjHL
Ee3GkHKnRWDlnVyF/zBLM8NiZ6uhDZ3Pb6/c1a3+/oNR9ciymMd4bgZ//4POMEC0C3f6P/KDIuGb
+dzbnSrOB49QXO3kW2jO7Lr6f1v26pitfayY5WkD0teL2k+Da6mSOa/fjqsGrRbm+pkVBz72Pid9
lptqXmlPS8k6Ef8OMp3uKVK/ow+Ze+jHVNQx4BSIAZfvOm8GnoXqKyMa3TV4/t/pMX9SWf/ddDVt
aFH45/IiFahcYo9eoyn7lujwc50Z9HX/HrR3IQFjQk3Yz0Idv5k4uucSPexvkKZE2APvcKvcBcpu
ML1WIng5dhKiH6cDOH0EOQ645iQ60Z9xHHwI9OM/wHUbjkOl1VyAEW34ivtlT9/WlU9O4eL2c2oa
asBPMUxWKym/VeJYTmtxxj8z0zTQ46nEZ+2/aWaKP5IphsZhzPPF/I5mACPA0YFuFKehUZ97Mx+F
YsEXI5GYM+qZRVIpGMcVcxTxfnQI3Vm1i3sVbVrIy6NB7Lw+rlzwr4r4RwYbrNaNBIUwMrDeECzY
s8jZ/ZbqfR9zkMA9p+Vvoi1wMGaRFtbLVhbO+tzFC1xtra+6lm8Wi7mJiYl+V1VTFZAaarBu42lW
q4qvnc3llBKZgH6emz8Bf5nxdGXWjUOpgsSBhUzsKICHZkwQKmm9DmntEJqasIcjrKUgztYyPypc
7vvvPxKEAh7jQkTZbqaHs1C1FuE7b15hGZj/QBRdnwMoQiU7/0SarsaaiT4DP1yyx8P6WesYci2K
UfzoND5oDqXCm6GI7BaRHWwK7oh7UhlxoIOhZeH6fZg0Q5oKZGB+QbIIqW3L36sEVl0g815t4Or3
pKrIjxnS00bECgroK3okFcq97J0hLNYxmJBgsapLpkdfA+DVucv/7FrObq7icaqaPnP0ClDvli2i
lmDHj/gIEE6J39S/jgm4yxjRBO+6S+u6i80lWHGCTCVGRmrnxhVuXwS8z56ZgSvWq6NeC/puoMQw
F2DCt4Rp2j/XnS39c/rB8NNC8T03Wdcj0VAHGIXdY+MEuDWD3EjwlUFpLtmZqLNeT+F1gV7Gj/Ky
gjLoieAmlkomkTxDIXw6WhWRyTxbLzTbRjo+OKmtjPixGgbGGNfECEioC5H8x4YCEM5VLf5bKKK5
Fvw0Ggrd/iy2ga/LoXA46p4yWokFn+v2hk/ipkKsjb5pdWk77c/+GzJ+1B1OzZq+vtPt61EkuVG5
UXN6FUQSEfWYu8GWSPS631pbK+ss6rQc/VE8nInJ+cct+rPWxZhqFbtYqTdrVLJay+TQ13UhtbXT
SSaedpJKcbkv4reExr6zj1OMx81sFSBXLmkFDTaaZfSjS4gg+a6YbdciOrvO48PpYrMLAGDGbZY2
L3lAS+HsQivha4xlkHhdSwpfw7ZTfnEt4ejfs++z8iFJlY2cuTqVuaStXCgzRfnErQiPocFJ7jz5
V18+e/71BWsHJ9cbAbkl85xBuQvmzVaLWk8vU8rIhGYRZLH8GjKfmF78isDkoByhyhe+7EYic1Ii
iAS+VcLLpwQqpirs4Jdk/xTDSrfLFo3wkzb7zRQXpNPSoHpZ9tSojmKOMPc6aQRtpb+kFke6fDvy
SLXhki/0X3Lfc+5q4Mq6ULGkkVmJN9auIL+g4H6pz9bZdFvLkDlgJUl+gYUmaFEgdLCFKlzq6Qs4
qx6xjzfDjwdD1h4nFhSGhKUUwqpClRKQHs0qdMW35f20c4x43rPj1hUEq+dw0cggB0zTcLkZ2VgZ
MnxUTxNi5uo/hJSKhhoLWWoI74pSRYKglykVYsMBvYZUrv3gifJMlWce0a9wykDuWmpTchrP3NfN
Aftx2NiEeSIgrneRmZMARD4CY2wYiFyKyozIU7yyTAlEnCWRkT3KgLfNxXfRauhc02vpabLmrWs7
FFO65mhltI1aRZgnr5IoUi1FNVi1K2QFiysTCsjNxEehFnv0arBZTgwhCkVhy65ovF306htG2Q0M
fcF+8GqAJ+hlYtpsSXVYPf3a8IzkmmDDV9v9wbZZGPdZgq05R6z3vzzpMwHB7j6HYYlJ2p+1pcwq
uU1Zp4ZWusgkrTJnZ7mEBj+UuohEBzIk51Ac2njsnLUbpxw2jW1cahoPHaLvaka2NGY4w3rSJY/Z
tIds5IGZVZYJZ6grtIvek36psshQBmM2/fTCYe4AdO0W2qHvBkLtObpndmeqJ9iEFqf4Slqdp/9l
8GrY+wMu1HIf8NZuzNXKQZzr+GN2FD9WVNia8+X2zXEBw1RGbE55vFzkR0ta7aljdVNzfj+9vJO8
jlaMkxJcXGQt7w4T0sKQg1GX1SQwb44k3HG0zy/BmzNhQy6Leuz05TIbSMc2R3eAzjKCf6JPmPTM
9swcQ2B85urrKTYSKwSNfaglvbJFJCfJLjRP8vTC5qu9EoJD2XSgLxLO6F3GUUqPB+vmY8DdEfkr
oeGt+ORyi140pi7GlQdY4ktTj7LrxjCQ80nSNWvuJ3gdlrl9jtdR3gTLHyd6vPUXlwdVrqT8G640
YSUXVEpdZFrkQgV5UATEVIb5jj1G7OUQkNGvjUNbNs4cnGfqNq9iLNfmpzij9MUtMxEjO632RxJe
VBIWZX7sMN9aJEQ0K3QtMyseITDlebUe1ezUiYPnPQpd3uR5dm3NuVac0rv/Kwdyu2pX7pvII3iP
6tN43G7sRokHa+7b60UbltGpcWE+qCChcWPMWw+OdGBlk9SMIAClfyE6FWp5wTGepMbb3N0nGq8q
tkNIQeOBtu5y2teadGrQtl8NxIQ9cfIi4E+e6xV/lnbi7UIJiPm85sVz4T9HIMEq70S0bU2BSYPg
YOfgWjp/2cbAULRrD8iaPgHjFmfAlW4FtxiC7GJkvMrd1mVbI50x9SQFaOIFPoJP9CtS/yJuafvu
4W98xxUAMWK5m7ZTd/3LcOCWeQxCtmusK3eFMRBQDOhh/LfeC875eonP9ey4AL1DKEcNwgQiK5nZ
zup5zp/uuDjQ1KWfSDw76Amq6Uzmc5c+GNM2Emv3U3WpxgicXy1B900N2xy4FIDr54jB+uPo7dc5
x6gsOM8q5df1Yi56xdPh2XHKcQ9Ui0/9OnufC0CGXlIsE/WoAz9azr5Zx2j5igERT2Ed6i3XgQo7
E4CsKKxm7O2vruuK2YkYWt+4DO3BQ1ltGk31GwkmPHkqlsb3RzTqb5H0WycrgPdPVsSTkxIPEU35
tFoBbQlhkdOVevIPDmK75JUEtjAZovw2nID2AQlpOymZjOzWkse9MKvne9v7xyeoQn++dMIkt547
1HJ3KpYlIF/2iH/P+OlHIm5n2m1FKt22vR42ZWEMNgUMXfHJkAldX5fUGPI68nr/pwxmsxqpjK57
3Ll7BwzzreyOIGYXE0LVxhvxO0nyMCPxxda2MoA2chy12iqpW17cqKYo7yriAu00ZhnRN5nvEQlG
YOy7v5C1WcmVNxsK8hZIQub4EdpuMnl8D264+S8JIEFxp9J3FsmLjsOK4kBdfexvOaSQsUsSOUoh
BhEf4YMs3fBH1f3H9QtyykEYrrFDbrOIkNWxNOv3K1DRyXX929xgkeKJ0GHSu+8/Q73nYKfty9Jx
4H+M2uKr9WqRcQmBlYNO0psEZ52CTiMMrRmJdeOig71nXHYfOUJoRv2fObD/Bt7eWedd5SKHz2PW
Hga25SthD9c3CLTB+k2GYIjRzmvimGyhM7Le50hCk7cLXuF3AfQRMUnMK4clBg/iGkEh2nJMYfmp
q6VB8nBR6ubUUhxEDcg2bqQLzY0bgpFjmrdaTArGzHErPmkt4CHPCyCQ/4yVEw//nZbSzG+pAo5h
eVuGt4u3b5nLWs0g1WLNdYFbIz89BvizzAvRVTGTySDxwZDLQhhqDv/Wg0DAcKOXUVOOjQfA7OIq
mOQaZi3LTFHz+n/J+hlvChgkGb+eQPm3VMqoWToZqabzJdgKM0nOC531LFimfCpwosKQohmfZxXw
0u7q9Oxi1BqS6XLDtSFvEqrAbvWQDE5aQk7HTx2XlhXRPeNv5hM5unCdY9LvW4rLC19JDtXmc8AL
PP1dElvMGZzhG4lobblh1vTvziM+U4aKAZ1XzFtGUxqD66AGFfm6mZBF+6Rus3CLNWQSexBCEsoV
2IPR1I/kwewNtwSD4O0AowzOA7NH/D0CBEBJuOHL47BW9KJKMm1sVnYq3sPj9pwzI7liUYgnlCmI
/t7AL/bPKCcax8tZjgV5FScQwCawPLdmJmwFSDsTepmlU3kx1ASfvbc/RUy7ikb52Lmc1PJERlk3
bOJP9QkvrbjhewqLCTi5ZRwL0N3FUSDdINlG+IN8dT7Casj/sxDg7rjubvRTmVlmiTncW8m3zWRW
IywcAIABxMCI6cBMMSiPRNaLMvmocOk98v65NJceW20B0gs2fBun06APHE4byps7Pzq3OVabBYH1
K6qqFhsPLdm3Y1hI4aI0dn7MKTuhW4EuEjQJqMdaafwve9OntWzM3QTk4h4m/lzYVqN6CdEsFkbp
pPdqkFixcvGOpcAuN6Yg8mUXir7mq0UUmwB9hcQOqHG5qZUlP05bDr6WZLU2wh7ljMGSrT8vNOZi
54z9BgNKbm3uEpSihEeUAJ7sog3FYqGpEOhRyOF8rJlUKnsNCmMv6E5rdX6Kj6vbPvu/x2WYb+Fd
Vjq75Wh10gY8Eo5YaNoIQ5cFycWBaOexTALRyZZ186ZChvgPvQ/Fw3w3gU0DqXfYHh1xfTkowVHV
cE74Um1ge1xAIQcGdWrziGcFpyI7qDeuVi7Laf7vjyiEMx5/4GE7SLCt1RpeRl/RVX8w3qTgx8AM
k0b0F+wKpxIRuAkT75eLhhWAmx/tkcFpngbECmPcDrOGqRYkMetAIHndds6WHFk03t/0nkfM8PAl
7weJWwc3vj90nvOM5nCzA+tGlm0q/0vEocu0I+eVs9MyaBnSMK7wcZrljQv+8qb2IwqslDQxXdko
5oEaEJZt3pZeT33CEzPOPimv0UvfMWU5Z9nkWEv8A7iRI6YV3QYv8ruZ/uRxFyvykoJ8FDyG7JC5
HjXP29Yj8mJz0Pf+PbH0rCE6btNuSOJbDMJi1cpjZMnJYZlx62p8gt8c3vUwtzcluIZbg337CjZN
tVHD5Y+3yysaPwTI5DCNU+aU9ZRp28qjMc9LpJI48OvNGvoLf1Ww/xzzs+oRpVHWfqFkMnuKanQy
sojskb6rWGbFZbc1bwJVPBGwBKYIAxM6qXvxcIXmB1tjSp2j1l0lZXCQbwaRCr/PTQpP8q9RBqSz
PPIAPa13wR4H+Bb1cWYqFZz38jKB5BxWTsNqbt5eiGCDvCYnlXdffPvUNf7E6+cF8n91cfjeznf6
QXXoOnl/b8TuSNSMC9LU9KzCeDPhDhT0h0A0UitMas26DnSvnNXc292D4ghOJ3+D0JpUl3KXhUt8
DKCUksUjUKAaldoMOtOkjMfDthIKKExUudAnY5Kza1/0yeTeBTKfCaQmY50FfBMJ2KJXqK4yYezY
+Fs353E9yFGhj7jklX2+r8iJmtbwt+RZ0OtbeiAw19j6O3yTXN5iotRYKdWqCjWYMLu/NIK3G9DW
ZswrBJrfk/LP5VvI8wHPCH0/jA27NpMFrUuYz+5vk4yLZiafKcPYcZpb7BWpejgwzxUn1RCge7eb
9Pe/CJIJVY9/MoTX8WwJIHsdOuad5wbGk9yblyenUtY7ZyEQNvWfhKGISfnvP4/0+/012M239N94
uKFHWaToGkrCodUsSGxZBAWCBVGEdKIPge/SP+VPkSHf7aAz8l2dHx9osK9IcY3hfp9OnjNs/duH
liyJkO5Ntrt/4B4x5TyPlrhWp8H+PkxSIl++7AzEYzZbM96cTrOqz0NXma18/Es7kIGMAtHaVtzM
I4Txu2p/5nuOIjk1HV9p42a8GTd+DtF7o5cDLwzC5VEE/EtWeqoEd2KC1ERAEVz2Py9enaKs1cFR
N0uyqQy0Q0kGoFOP7Dvo4dyrzzo2BZKtH+2TnWtc/ktagrpnmayogQYa625jmZiPOx17EV5hlZiN
yFQBrMv8AawbmCUtHkbpkJKMTfWSdX29mNs1/rfwTtKIm9HtoJhXbCKCwzRAuTitYImhas9752DX
8NPpTGhTc2gIIGCBziIHKeLluk/9W4BNSIPt5cwnIcoWE4er9QNArbOE1dLGesZoI5vKO52EkQ/Z
2ypC6B0f0eh9ZH+NGy/2zE5gCVUyXjci+JWmX21dCJqeZKr3UEvwz1q3FSlWz12SLzx2FkK1kzUJ
wGnaKt23ofsjq2TT54xTUgpriP6nabikZoJGVe17/HhMopx3yeIXCX9TpYbta1vvu44tVFOcT1yf
/xl5TgsexjGJ1p6oTvUiFCmYnoao97d4Ocj1CtC04+TUTbKFQqtwxAPKZ84LPK/QPur8x2PwlT5i
AwKH2RiUJo15OCFKemtea8EqbOBGS0b4H/FgErhX/amS+Jn75fmoN5mvHum4Qe5TdURMg24eg1Ai
QUC7dzpl8UsdEwcZqUPlxc++1+t4LVaThLlNRvmQtWtGh35ked5CIipKZqb8ZLxdf6rFrVKmvFLO
Za6ub3O3c4wo+sIUp9R5LtqXJXoBXO6/bneADTLCZqvxMeUuNTGKW7Un5boNTxn6hOsoHk4DxYfR
q7+PNDTocb7E3W394cRfsrE2XldRNAh7GRRai8Qs8eCjCjCDoZq643sSJhAeK0TdVNHLRaa3TMm7
SXM+6wThFldS4zr+DxxjoP0sag/uoBtGhx0OMi6gtmZAVrQmEo+kwC7u1vMeVrF3C1xngaDf2p2T
auzcvagxvRvccWqMHO8uN0x0FH87iQap+ibFUn9gGeCPgv+bvrmw0P+qR81xgMunJ1sAiBtxRRFR
76W6kAZNmFcQIBdRLrs45FeFXfoWR/Rdu7vy7WMoCB68dSA+MRlzDbTl9Mfd4ytQMAn4y+vtgoGN
CdpVA3tTfg24Z7muJGrCIQACnYKNPbZ0rCZ5xbWflLHip7qe6Mc3HJLm7qHGch25WrKn06dEN+8q
957N8wDPlksxvXex+vqarIkakXHwtSOpM8MG9VY85/r+P/TFoTwvK5KqZID61uY5/K/feDh5aqt+
WHux3DUYQAUVWCsFCmRoEuhCi5CBk98cOaX6hc4EE9dDpXH+EhjzimckG3T6sXv0SXPvW2TIqrCM
PJUMo/kbmKxMgUGI2QEssgH6d+r/rNBJEsT2u8iFUGG0hC5Ri3WvXJpEaADGWHyvj0os+gMNL02A
aJ/eQpTtrmEyI+zfzQ8yzuSgRcK2d9p4SVkxF91vVBL19NiLnTTjNVIBKSpxFf4bl3VXcBC1q7e7
hrVn78i3hT537VVR1Gp3WVcqrUVDAtOAryWQlIEvXf/N4bMqoVsQfi17UNfDO0i1nop0ZFJ8R7q1
8LE6URFR/ZFDztA+EQFC4lX5NZAq4xNbJReBeLU3ea56BK6qJDBuFqG4XpKSQpMA0it3mLHGA32q
PlIuJ4HdGlWLxtSWfx4E0mPXmLT1prCZSdQEGoTrn0NM6DezQ8JuylWkCPXaZQOtSB9kH7nzvM9w
L/Fu8JYKSovObLWvANAAT2NJWS63Qrnh+O8fT6GyBe7FOoWgern530LpcS9I7jaHWS7Zlbo7iCs3
+wB2h+j/vloWn5Bab6rmiOi+HUI184P4pH2vmNYlsaft113iALRFs5azP9qy0CPktCaOzJbNrJAj
AuDHzvqIQEYbYZyi2pzOKf5yUeuJ/FEmUhR3xRNpsHqmx1bbvx3brQirXM22wVmqXs1SPxrNsot6
PaX+GbyQmgoEjSCtPzoJtfUfvf3ZQBybheXhWDdgZcoW3zfQhNV86b7chmLWcT3nUNlvZ6ceCizR
ArhVDZCI1585JjGNBxCBI85Ld0W/I2dDihD/3UzwlYtN9H/LAWOwxGLUmigI5Zl9tK+oVCFK4m5+
C+hi5osvYKKD+FL/JgGNyMtal8moiYQIfmG0sVZuJ6I2IV0xdNqiJXsTbLfhbxwb7bYE2fAys4uS
Yq2ZJYEkosgwzrNoipDx3VFOAsSe46d7KGL6K8ToOxGprRksb9wML0yBg+JxXbzeMCcEjQ/3orRS
c156U/kVT52wbNtuxoYzZiYfjrlrhcajaAP2vONxq7tuaOhiWuwx+WhddYT9wHv0qJKA1ZWq8Ky5
rkOjuQo0TEUlfK7N2l6rGLTh6t65lo5aEaBQBL1mu/IgPEx0o6NC+CN5WJLjxRdCZgIsrdIEZjq7
JTPByLGA76ao1iMiAuOxTter7ZAfinR1da7mZBsOqqf/dEJy8mPx2HZJSDSc7MEg8bsoAYZ60V/l
WZYB9iqx2nc/fyDCJUCYT6RXCHMT9/mOabccDHvm1CS6Mv/AejrxwvC98ZqwUUifRl4SVPg/y87k
nkaOq+ElzBs08N1ZyZnNwzEBj5Kx2/jxBCFUqwx1i67PYvlwRH0Ph9fleFbpQEZsf942hJ1tHWXG
XHoFWrUKoccYY4inBa8QNHRVdARW38rZZrvd09IX6OBDSvkgAym0qb1Z4V0WZwW+zq8AaoR6NCGl
AnYTKw6oml1iciP2MEpjo9Gm0YEsvvnnvTbwq+EW+0+rvZGCAJoAe0i1SwNwVyqJUdjlb1q/mB+W
9mjWfP9aUBFrDXEMiA/Kq7wq105wyX3VccsBJDAHUdN1m0PeenQ4XaWfUbvtg7LnnN8oSSWux5UR
G+GQ4VSX2wNf7exV+B6EZRwe2gledQCGlFsqwXAIz2u8yJwkzvZYtTnRJxpo9cP4CIkS+nMYpbcL
Ehzn3Sr9H3q4/ntYF+dm7Eejy1qYGuoNQJmQSP9YPL720ca0oI1KqZA4aop9DWM+N5JQkUG02yMz
UUUTqJXwR8jIeUh2BXBnSzlOQGg9Pba/QENjXtzRzUmg26tYC+7R0ISNI40o5AT+ST2r0HvgL2AP
nMI8A02V61iKQU/a7MW+xcKR1xGUPyuIRQsvLnNdd0qUHSzJyFVuOOe6D4HBTcB63OOsJ8JBAyRc
9sYWDh5nb0mI2Uq3IEuyI8bh/nlH1yl6HfP7RX5cbM1Cy6r/AAnk/dAIOQnJ+M0SQ3vxZHZuPHdO
9P/CBdvvlMk40vOumitvuXP9ZCS3E+j+riB3oNk/wFRHwznQUFufesBYgQgEY8X41SrliG4rmFoo
0hOJatG600dYmGABBV4xR+OW/SrdZ2sK8aRQuG8BvRv/G0tQ7r57wuvYsjP9/psvoctLXXHhFYZY
9JfNnCpbOkBbDzCI1LRvsf2Z3Z0LR1bOkEnL2uVhrfocq2h+CEyIGFrZUf6Y2wSMz6ArHe6JJqUZ
Pe6oZ/A5+zglvvL21kluHB5Jf5DNsVN5N8ysz2dMFpQF7sZ5bk0Z+dHNjPwr49AcuCRn/Zf5Kjto
v4Wt6vEf0q86KKcIVRQg8wCcCf/5MeHm4tRCO0nmoA43625Wtz5sv4xaZDcseI6SIkTXsusfbiEN
HoEbgoF2A1yPgmmZuinonMDcqAKHbGAyYvmGRrrTFPRn+QztcwB6GN2+Cqj8R8+9S97I/S5cHjGh
WvlIRf3FtSfSgAbogRS87oejzTjWCCIeVpfpkkP+its2XqQ2Hmrj3gNIWwuGDDOjVov9Tke8bHNU
eUHAYzn4vI62SAU65OXq/Pq6AatzU6kOX30XoZS12XxJCQI3CNy1/EoWlDA2QIp8vJX54X4Gl0Gk
SWKsolNgRmeZ8SHrtysuXGSUY7iDWae1a2X4Go68S3AKi+CgEwzPTGHHQ+6hgxzp4pa/RpNg/1/3
v61tZykaZXn0eLdD18JpfdHM5rlwPYES4ZjsbEWw5v5spUdKuNuaIRaHKKLnpdjTgoeP3ZjhvjMm
YIcvByunwdjM69U3KNlxc35363erlvS71Zmj/8Q+KzU55CHmw3qX6DhBdjTEtuhIV2+BI4CwMAyh
Ds0CKLvJX5bj2ucTudertQH0W5Rh8bV5ZLCdCN/wC6mpmYXs+/yCmGCnjtccayP3FYPHHW4cfZNL
Jr0d7h1lQwb4YhoPcPjaDSRjUZ4R6uR/g/zsnp4uCzmwSDVcpPzjVcjjog3Z2+4xrnhH923Uk7PU
2jHsx/nw3etwt/cZgG35jsrQcO4BRMu5PITh1TXDKJ4P6W9OuI4DaMqv5p6cS3xNM66FdiCr5Cb1
/7gZsaqSEHHN+oLsxnEizKiyF/R7sIwbZc43BQOK5uxVOEibP6oXfc9yjGyIHXccUwavBER8aSgC
CHbO4uWBKmL4oe14dAzH3iG+ayzFEs90ek7PekH0CI8PWnWHrbsvMJ68s2CKnCDM4eVmk1mtgdTf
9Nj7JOGMwmMps+GvrTpXKgO2SR4zNFHjZRKMYWjp3ZOqzV2IirN2YJHHYtaoTYZ8bPl6LUFEH+7U
3tR5XbvQ5HIr5qh1jJvDxS0BnvxQbiQLqx696skpMkYDIZnPfk7QNas13nvqKNgrBUVm91LLrqSO
Pfu3LnWfy0yxSQ8exx3elI4v7OWmf5mlA2sC8BjdoIEkl7nZWFc6nYEEgjnewopp08xMLahD9dhP
MSzjRKDXzB9AEwibm1iMYsR22wEDUU8RnhoRGiNRrrkLoeHu+W6fE8PxzDlbCCzopYo5j97GsEN+
5YxxtYgFWRoUm53FZ+y2nOegy3DB6JNTxpC8kGv2raQw/p2s4iO3GIbVmseVo9O5Byn48ZfhzwXY
jGg+1ih940rhKBReFxamNyR1JhwFifgIGqtUsk/x6ztOQcRbOqUkiKyE/tKqCVs3djAxNbEU8SiS
D/5bcH9+44DFyH+M+EFM67goSVsaSYhrU+hDUVBuOSSwF6XTYVn8zcq1wNhssiK0DO44nLEHwX6P
jAx6qK5I0CLKHrUcCz+f4/nP8Fkd1+mR+cuz8CeEeI9nv8KBU1/8mKu57wmUX3HZ9nFvA29cp9ff
x44NGXBAfH3ANjIdziTk45wOtdaVrTJ5dgFBBmv3K5nURv8kJYC7S7x4OZ+jOsy7bHV+Uw19zh0Q
+jd8kO8+yI7CCJKptp/TCtyaSaAqigqQ2OrLgK6rmBJmcLZbO+ZU+zMGN0oD9P1q4EBnPgRmG0JA
za70uJefQWtm+SHU0MgwPSVJfkOjOPBE45X3bN0v5/vQEWyaIqycVnSRZBXRD7XnOayQHVATZQqm
+o/EzWnG94v2odOxtXCk69qnayhb6PZlkYwsn+vawyFrx4hryBZhvuD57TEyASq8Turl5j5K50GW
ykpoDZc0tprqXsQ1CE9jVE4PUSmVacI5r+6XBYp8v8sE2pCFgf3NjOlof0bvAK8pqXT+TV9gFYhw
xEyPoXTtN0TFQ3rbpY9V8IZ+hctpE/gZzutOewai9qv0GUFr0aSA9WYuDbjuRbytTtufTNHfHzIM
RHPPFVtMHbT6piDFIp9dLviqSB/D/ogbxWAPKaNcCmGl8OEGI/KZcEMfr1PPw5Vu5Ta1xGzYgnRL
22o0R7E3S+iraGRmLcI1UtnMKChZH4Jf7WbPRRP5SHaL/NS4ro/STk2CFJnqyOv2BGlVi/iPBf+Q
yZW1+1SOBZoc70MrsNw8f+sONFx8qzNcetk0+yYou0m7EzNjAs9XQK+rPBHSH964oNDV7JubhFsY
9NSrcn15+zEOZFUCBcV65/y5+6LHGMBjs5VRu+Qc/GR5j3zDO/V3naNsUG42b9i4T7BGactpKOue
KlMXTsaAbCZ76CM+LmoDxoZ4T7ZSuQo5HORZv5m35ff7mhbER7Ka9Jiivvhg2G+6U5fFTWSwUVvu
8m1nhX+XCt01fOJ6G9uEGd+9QPfS9IvEjBmbSQ49WB2wHPQNRl7fzVy9ltHTcuNX34BCrBHundQa
/s2oxfKAm8WO45FFnWGUw264Te3e8IrK+eF0JG6AErbAph/o1FSNmykavax8pM/4sSbc6pXctpBv
BOyokMZsAcR0yRilRABuEDyxG+scQV22vFJzbTEjDJc7S2rZKfsqalhEJS61xDopec61SrXqsR63
NWlGBghUGnjAGehuVD1uLl83g8lwQCAbFL7ias0VLCV6IMx3xx4BFvv7GsSB75xpxwSWm+nbnt3/
REb5KSODzT3x++ZLGB71Shpt452eoV/dAo2sxxgqWfQqOnqU3vZZhkzd9TkVewF2b8mcfC542NFX
paj8/hYsGR19K5F4Ii30NvhoDiWgntppA7EwOWPoUt+R+/xSd299KU8vC8A/exc2qQwy+IHh3/0P
704DvcG9iH1S2+V61HHtvRl+4b7pLFDjmQkUgM5UpaY8a4VyfT1OgT6aVMnM7w7+ggzcfyI/qmkH
fpPeaoWD1Zqm8UFeebbAm3kT30htKSMsHkRem2+NMOgwFSBMZHHxmTidRv+pBrQCEmwqvIywTSO5
gNwBrSek5OR1luzT/gq7ByaSKsnq+3XvKsOThLfn1Ex40gUCQLLEct3sgodjqJjhzEgAc1avZylh
O2wHKmY9KxCNWHaxIBQymcCuz99eSvasWjZfLrj9BEPcmepEHNqoQzjZUf3UZxyP9zB+aEEdcTsX
byiV68aP4mT/AKGnfp42rzG8ussyve271iEI7eAd6GTPmDk69J3xQQX3uKZM+nqOqS36fRgqQZDr
h0VC27aNAEZsDJYY7a3B0oYVFNC7lZWMfJ6xBgbc0PHaxnHfMwlVlOBidrlAZRHXM7nMyzs3AAsP
L1FJn8ctcssL8uJiY6IqMpxnG/OloAWfynMt85iec67vWPA9qLIiEsKk9BOtKFTPXAcKleO7aUxr
+deTUjU/SqtUu8RTu2rGbLileA0D8QhYNS22fxvrQSd++cjuKRJXpx6t54N3VJt/b/2mpXw1QQ+6
CqVioCHU6mSgMP112Vqo40+t5JmEc2y00HFCn4pkqUShs7s5NMq95bh9hy4ZswJ4XkrijMJ36/OD
q/H0nEDjrn7HU7Mbo2yRmMMsElQhgCt0+9mOTmwPgUhQ0cJR7EYfVpK82wINv5hBLO47t+OgFSQo
hw0v+27D1e0yYMJfcEJqVlIBZkR5vUDlngNjBCvT9igps3H3d8M8SF+UElxEgVQXf3nxZoDKih9M
UgCYkluqExCSrk6GQWaeoehzEhmT6tJCiVgjPWEPBoPHFJdtyYYaXbv3yi0HPO7bRJ13x7KS2zIi
StLAQ31a4CRNr9szPDuBWpqhaim2iazOEqu65JKGXcvvvHRrixQgbt2aepY0lsIDOqU1vadaDa47
swzw9lmBJSMjNG+odozGe+S5Cdvr7B+qsCbQY4mt5lZr9ywLcQQz0rgZk0Hnd/1ghH70T6GhlaVC
2A7IXuaE3aRhpjI4vB2yJaVPIlj6QGcakIcsbxUGx0b/N/FX3EiLBQM9alDTUEeVRh5i/sHh6Lbf
2c2z+oXst/T0M9lmHVpRys0x2dZm/98HyK534PLS6Y8nQwLDaZ+erPvpeoMEC+b/IZelXqdr65OO
fB/Rwz9K7daQh0nkYo92p7vcjd3P48lLahSQWYH19rDGq7UelBB5H5F8UabDpXxR7FaA9XdILpK0
y824z0f/uFGCkPWQCOZsoWvRCdp2pEe57+1X5P5QxhEmRpOjbsNyLb8Gc3J+hLvFYS20C5yG21IC
RRQW0zHaETYaw4921/tr27UG6MsVPNvRwu/hL/CB7rExKcPe0VieQpDcye9fgq5wV5dDFbYiFlCV
GKOwPPEHlPkHmuvyn7TkwkAKaCPTJErnUl1RkCFey2ENHhT5lL0IHgdjR/V2Nnua3Vm2Q5BZIZ7e
weBBxiZM4pqDSJLooW6b6Lub3MBLTcGaHS2Z6+IRGSCCemD+vqOzOBTjsPsY4aah7F6/C7EXJpEN
bhNqygScqGjZyzCqmPw9WXe7xkL0lCORzvJzT88mIaX2x+rBq5bcWFgd43UBfFN03oFPnQebSBnN
Mj7zYvb61iSlpYXhsdZbfNzqVDDrGUx1gUNWn+1rJ6wH+QbNHP9PmA7UUuPFkxXSQqMxgWCu0gOG
P2DKR5wtGue4J674kUCnCFDSyyu8jRByWuVVSyLqukZafg22miO3etMtMt2ynWtnwZrNPTTup+Mg
+FvrbKjyd0W0cqzkEhC2HFbIFeS9h8QdSXLADRljHzJz5O0HnqlKov0PBiM+arXLFrEouaKXAsWM
mr5EvKXEilnhBB/hjKLMK4zzf3+rZxeWeI4FIEVkPpUxGl5ju/UKycqGq4K1sgtT5xqbmZ+zQVAx
EGF+1MY7ex3ob72JqAfB3XoQdyrVEPGYmIrLLs4VzKSWUs6eKg5rSIRbMoh+VKsfPrnpk33wR7+1
QGEQKb6U6lkR/E02hH4WwdSLL0KPS+MaYHhKt+XPQZeZyzP2SCWmpozG1aKp2qlKyNPrKam6niSc
p9swhz3yAWOl+TtSMFsfQgJHbkUOF52Uywq+kNnLbsXcC7EnPBK4RgXn22KtyrAfyZBOpTvZ3+kX
tGj4Aq8oZKESfqs/S9xK/jnFKCmfzsqCGppiIhSXFJtsSQyTtX6PRcxxYu/L+3J6FvI/UGb+VQe/
rlIe1c6d1vzO1W+cODCNlptYvB9deSbd/Vu2kPrAyooMvALVSCn1/yOVcLz0VjHywmeV2Pf2hqsu
AwjyXhB4aPYAANd9/eqNuBuy1ywH9s/bxvqZRobr0Cq8qLoJ7trcSeUcEuqIlMm3QkRBXiFiYiTU
N681i8t60ce/fzzQtaBQmwlbRUdrv16SpbRzVB0azqmc1ydLId4T4iFAPIIAucjz/l/dHb56h6mP
vP4UOPKYCwJJ1b1QmJA68u88iuZpftLH0Ztb49KEZBa5q7D581UMmSPHhdxAOJJcBG8FF1daZ3tv
Cx848DvTUlJ+ppj+KpWC78RZjsU8XvkF2wlDR5KmNYezzqj9Mw1qkbNvdTjm32rRFZd/Q7ZrEyHO
QQop3tsj/n89e5pUCnSY4K9l7frBFjcNVYpoc4v39dbDX+Zua3blg9Kb6ycpZ/6ePw==
`protect end_protected
