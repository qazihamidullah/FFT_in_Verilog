-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
049cI2Z6BoHuOIbcbTMt8Qvv3gi/UVee5p2I7kNKaMUoUvjjYv09xQrf215KlTrI7siUo8tKQhJw
5GKPv6u2uBUl1FyZIsDcKmG/3g4Kwvc/SKp0ZVkc429pUzjZd7Vw8/sBVxf41+Di44TFrpTS0dtb
po1MCwR2rgMdj/RBNSgrhWyr4hozFxa75OHHAA/n085Wuz7+ByimSbOc41lxRxkcWbSOz1ozEHY8
/dN/YDczpfJfbZe4d+Gz2Hhk02Z6Qf8CmO15Mcqlm7Bp60a5GHjKgbUG5Qg7kiwz6CM5KzSESrWP
Ur3DCebPh9Ikq8jTq8xZSpa4/ShoQQsLlICvsg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17008)
`protect data_block
GlA+zjDYRqPY4ck0nyY7x7eBCW7QB9rBKoScDEH4nD2uUcXU/QuKDTkdy2WzABODJyGW0L75ixTf
Tv/es+D/NbaBtkP/ISJHD8HI15R6Rkscom1A1hc+SLontdYFg1jOn3s6rZykmmIgTzoCk2eQdEr1
Aa0x5Io2Gxo+rj4F7pbsXoicjKhExsbPx074W8FGsA4WOW3yRaCLPJqpsVaO+2zRutIXTczmQJPo
hwJ6MLwB6H8xVWDc4SsgWMeGKqWRst0hXXaEKH3dEYVkZCT4/xTm8SXSngMVHgGdJ3bKA9PvB3Ea
JAOX0eshELwAjgxT3xES97r9ks19+YlcJ2SwgGZjxZbKmJFLpQBHZMssvx99m/LGZ6fpQnGdeMRj
yyRxGUX7kBSAxnEDlySNFL5YWcfix26aq8qSLA6uwHYSp+vPVIxhPVOW3WH4zvySsan6/lyrN0X4
Mux9NGBtLOQrq4muCzWDpvuRBC/hh3tQy2Ud/gJ96MbsG78enrOqPYQ0pxlDw2G2UqoyYYvIihut
NSVl0KeVHygEl2TawZ+GJjtkrHly3asIDE6qNvQgacVyjH++FvWzjEcDs+C9O54cKKDnKG2EoVIX
57LT+rBzxw7l4HynNdUw9j/w2i7r8vqp56mL6klraev8NrwY5VDKsTYKmf+tDqqnBttd+eNGahKX
G1ubVXvA40Zr66XhzpDAl2R6EzWHXARFdiggi1zECbZ8Z3Tfg6wix7VZ6/f9kKtHas+p3VTyqSjA
t1VGkKlFpHFWtYTszRb+sGc+hn56UFKnEST4B8i3Rc8hJNJzh0yHwDAeMnLYd/5fYPsBCxfRbL2m
59WEKo5FfVTwpuXYjj6I4zqMl+qeLKuztU7o4AizWAsquck4U5fXGjj31S9TC6Q5AYijW810CxBf
0EaoeSwT1XnBCixB0YvYeOvXPWuduwdjyog86xoeXfQDvVE7g6YZfOL95eBI5JJeg2Fn3y4PDp1U
nwYBAkog3SpO9HPTOI5W0nwLlY7pi9H23BoICrifDhC9rqqmBQi+CFvEyzG6HLtlM1UZCV4Zpn6n
cMcih3nn0UrSCUjuXkanxA5M+1d47AbBU8kwNYAmzgkgSovppomSpyqkhhLqukXCr+3/l6CK1cyo
zitO/SrySQkhdLgQSQeZsKwmoakepCBXqX+7YjYdEwKe8xLJprLUiFdVd07M7PcmO8PIFPDmfEes
Aur91gDXAIad4t26XtoyGU83INt2Qubs2ffhypodEJ8o18M/2wBL01UtKlGZGiCzdIEKcXcaQKzF
9tqFwU0q6oquieFGzKJyouRkS0yNazgXDqk7p+CfyWIlP6oTavdeeOopVvYJffkv2IoqdTICN+tP
c04EihIxy8n5Gyysz2uM5Jtdkr+vRuc509r0hsXlwzcN3qHzX0scZuSuge7HasISeswkY5j7d1Q1
h1IpYSTcAhxdioMyUJRkAnHy9VDXW0MxG8QC8TsDXKTcxLhwfh4FIQgnR/IfN1bK21i60sr7Xg6w
q6KDe7rSzWsZbWy3gynDw6f+C4MpdTE8l9Y5V94fhzUpZOYlYN10/yPrKlLuSp6AJuHZlfaUrG/V
LCZgQSlLsvEh/bDFyxuCLGRF1pvyb2APDmOB1yH6TLbSyn6PkBBemaebFYiG6Mc3Ol2Npj1Kulof
jB5PcJfjmveAP0wTkH3b1seUSPe9rlCuUQTNzlbQnggXichsd6+fxBvzMG75iOL679A5Pg6GndpF
ntd+3C2lcT5FbarbP1cpTUpPUEXN9Q3Rdjw0+A70fEGedkQtw66VnYHXg/rvbhlTtgIvsYfrQ/se
7aoK8ST050a65YgnMAMwl4jpM/zyik0jWy77dIcRiH09XXenc1wuCeoc9+0SKCI5YrYJ01L5Hxex
PvK++EjkKM29OiF2NaKfX9ACPawmgc0xmog6wFupl9T6VUEAP2nNt4h2GvqxBGDp0fsCe8g9BXWU
xQOX1VOhgGky+urZ6EEtiZ5kaZrJ6AwtZ4qQ5PeWvGWTxTs8amvbENL4qAOuj4vjhXwRXuBHMR/Z
HnxMAsGiS5DqB4sILgenfhAoE44deT1V0yg+1lIIWN8RfQLE68oB+fzuJlGVG03+gJLU9EdCB/yP
WPN60vkd+cQ4ud6w8HMG/cKp/FjYp7MolalWJx0eMcaT9bXJGx4hW1jDtIMcSOC1xdNKCOVfjbDa
I8rF1jplgXWYlI/kKZNCHu2v1GZeSSau6r6ad8WSSW+qs8KZWKp0WrXeBcJYWHnmaQlrsp2uWskX
4oMpyP+rnsG7t00xtOgujUBVsyDFFGnYizOTdq04pdI34dLV76JFNZiEwfX6um0Y5JQwqyShittE
P+FxBdDPwPhKo3j3+OsaaNSlJUZeJGW+HglZ/tW/J0y2vo7k+EtokF5+6y0t7jlqGjg8YeUsnHjI
2LfSEU7qT8HZFFKdVGaVXXGgQ0gSTV8AcqnzQWf+HmchOwQbSOSw8yp0McGYUeeI5D1whozbf8Bc
MK459+wTN5BO+HXXpr8wSxhcNzBo5mjf5zuhRD7K92NPC6i/vUkREOG2NVIn4ez442zi1+H9fZLK
Sk+WoqfFaEfgc3hKARKiUg86V/59hajlVjhoJgLmo+T+DLz/bXI1eTfhXmGDGcdXeFaWchJf/Sm3
IVNxZrDEZJvZSrUWuR6Vqe18qPelbzPhIK+QWRuWTdmM6czcRLWEYDQ9zr3kJFWb03bAY0jvd05w
VUlhCmoFKmI/mny6fjgchVfTjN37Z8WGGPdOa/NiF5RvQv5dFhTPnxTpVuTfzxVOh6na9J34V5h7
n+Opfhu6Zm0+t+UoMBP/axpbNhDGpgoM9niO38nuyBHunXDAi7D7sj5D4xT1elK512uo8NKULJNc
Ctq3uYoJomjicX1fzZ8OSPqi9TDfXQmBZ2gG6bi9JhVEQGcPq0qC6pvNOO0Lo+z7mViUiqy26nbO
KzDKzEGBq31hXTrKnWzBXF4Mm82LVtKD+0pE/+cRriY5py5OkB6CU+Kif7KtqBfZdd1nutjhwP0R
xtUhbm1R8r2Fdr1SNSQzgwH36H2dqZI8FhWqrAS/+/7hrf37o0gNeOy5/irtdoZtS+uq2d0piRvz
Eu2sTyrMwnb8KTTxIAl+8O+3Zj3JQwxCLRV2hPwiNwKbRmt302FInMg0UWTSwNAA34HK8B+xPhId
LoBkCtMiCh6ZBHAlaaS7R+Ma3Z/7q1+eapYs25KUESPl2JbHviKFtGXg9OlDmevmHfnDD9vopMzX
f2N1bxQ2LtMPluNVu23rG5FBJoGD6gCx5qZ7ruP7Fhl1wDLTEGDY4KfZIbyiU94St2X+skHp9a9Y
dlxRWAj4ALfXx+DLyFhn1xKb6kM2buU1iuIpm/HxSnqymdXC01g/uiBXmLcHOniAfVfxfsdcJagL
UubYobybgxs0/Ihft/tZcubHT6dsA9gmu6K2i27KHQu37A5B+uorHO6Sx3lJxzopxkVrL/tpdLfM
KYlmln6JgVZG+humpcNhqMz4Z6WgXcQH2uYi+ayZlFwzQCqU6wXzTU83QEIvTePrsEopnKNbde+3
kOMsLTX6fp6sNQSD0uv6jUc/s+XDiP/L+827ef+2Y34mqJchIgD+SSzm2V9Ev2sKiIDETyNjaj41
/p8/Pw8qIejEVuwiyG5tnj8usUV6G0LoVKAQPxIBaxnit45A7YWsC6yJ9hdCnkuvHoix6sdou3Y6
tOEX0Py1pQ2LNP7bx0MhWxn+zRHvgeJ9FVAtrTc4oUBaV2RjIjMUEwq6Cu+PVMJiCgLV1x226y/U
+MuUJC56mpr/Hao9xCmqRw41XLOWfv2rVWSq1V4oqDbWIKd+Mb+r97V6Ye5qlcuOBp88Eu+ok8sc
iehvfXVAn+uEUQ2AtIR7zrxjGeSNDanbk2/+t7zmEGup8NuxcWCakbxUnnJDHk/0e+xOGL8n6OhG
BMpcJkTA8Rq5bGOV5qjniYBMPTGHzRiWjlhphNOWRIJXoAiWUS03h+deSNjphxsQKsEC8W3Kl3IN
u+UQL7Ku3+d8b0BVOn8PeOgzmyRQr+8ywNEgx81Ju58dHUifW6kYBYXSwFpXb6Nvi91iFAOTDTad
JYPjMiaHx8p7Z4K2kQ9yfJRk9ZMDBqI7Z4wb2cwaU91od+17lgKnn8tN3dtva7zKW1g905HidL9B
Zskooh1G2Ku2vcpnzQSI/qDy05Keho1jSHsegTeNdTdM8l5GSz2ChZwgSCg/xc/nG6ZCziyQL+Q6
yQDNRucjboN+1wdkJI/MgBbwQiSoMSPgpduaZ/2D19MLiw1W0z+9YDexB0uIfn2HPuGsBlymPD+X
pqOY128gNCF4qUxkw/1/4wtlGba0j9ag72CtF9jFqy22xMsoCIjy8WlXldBm+NE4E443lp41g2mJ
LW5flUqJXLbkJfz3fVH2IS9svzgEccoPQ35C+mZJ4pmbOubqUvwl8PWo9pRn2VeqROZQkxd5zlXk
y5Fvty4VQRt4UWFeG3Begz/1LtD62oQZDq654SYpGk81tqzKkCdZu1p/7x+K1cvdqaHGLs+9GVlp
uZgkwYKSvxpJyYoJ0MsqPcGxBFUZnJK1jsgrC2EcuWd88PS4s6cnYVf6QtkD7Ib/Of2j0k/E7sQl
u8rnMM0VRWbqIF/AW0nI3dNqcftcAbPGx6FvgKFZSrulzd+YcCqxmqx859ABohKKO59mbAl6+bTW
pWFkYakcF9/frrq28woWLubwv9Pdqh0ST8Ixzzseqn249gKQ6JjU5fzCwscW8kgK7ru6B/zBA43l
woNXMiMjLslIw/+H1FMQ9yY+agek34wKr7AXeFzsjB1RWI9UrLsW9Zx+MqG6PjffRJhewecOVB3Y
GVfJD9cYTdcfUZ1zYQlp6tCLwEKZfx00oqUkSzQLRYSuNxBPn58EeV5S2KyebF29YSavfNWUFp4n
7JNYhrBZKH2NOAKWYYA/H4tfGjunGZiMHiqVRIBFfJ1Vase9iAc1YVdyurBWg46f8CixHtncyJVF
9QNR0d1WMHuBNOOkVbjerJWvQphSss1LLaEP38XBQZfF2SQJFNtwOnGAZ0D0nrtCFsLaWcSPE4P6
WlKaZo7B5F67SuJfwDMWAvDAEC7Mj0ktM4uyGvJKqy03toIuLJ0YevgNhMOU/rRcQNo70lhIuAO4
WUiJzdl1RHUcPwtf1y1wZi5xXl+5h+SM391uYSxvQz+0g2GviMOQgEcrDkrEpCw6mLldchk1fCmO
7qDIpZVCYHkgABtFieOfDcfWVDLAl4p6zjINty7QprJbXFVWc1ijYs0BK7tafOgiaNoohhgQ/tcp
IykDEu6Y7ftgLOYtmBSlzbGeamYahbHfnUUlGi7sene8h4fJd9iGGqW1ckHELUlo8xqLq2CR+jSl
mAD2MMRPyesPz6jmpD5XzU77BU/co3ZHVLEjP9bhIOjQ+oEgh40HPdODvVbKOk7EV57B3/I+Zpio
SD3VSmFg3JbxCPJxsXIVXvO1e+VOyfoeHQk3idzQ2S60mezsQI0KnX3Jc/ANoHlPo7Vs+lsHT5Xs
cC7vaByD+k9iZ4xrpwvqTOX4nV1LafdlR7G6P6s0asjRUyKYkrshP6Oum10iuJBqsHfRxZ/3Oj7q
ONMm62dDm8myTKumrLbXxhgot6oMrmGazbR6e9YJgsSpkhJFeielgdV5wuYv1YQSIK+7UbNzIbuI
hnWl+/JSbMP1rF+QgjT6tjn1E554p5omKvHZ4bZXJU8JNo6PRmWM9PkZdp+npMKIh7t1Pu8zlcSO
HXEBcO5d+FfrjC4O9Ps4Xa6ZOVS9ewv4p4KooazALKw1EmMYXdudqxF8y8Gzt6bp82LM4pWTOry2
2AjTtwIasxO0SYp5lXBg4CJ6EXB8Nz7N669ztTk/tN9OEkmxTiSmFc2Bmg+wB/HvVLKpW+VDK3Ad
Wl0YMe+GVoYhR8d9ZgqM3Vd3OFyCutvNqagF0r14AvONE7RmR61ZxeNIB9Qm73eB9U/MUYTDogKk
+j/sxEnpYIN/Dl6kW+OKmJ/0Wu1i/7hqlhVcAb+OQsmlnTinb73b4mJNKhIsp4iqT7Wub30e/NEf
y20Adm+zj7ViZGIna+TKojctBNc8czhmYuWE7tA4vVw+u7JwSg+KVfdQ1gHbrHTZdmuXPStTPoz2
WfDYJI3jJd7x7+NElsnVtrTCy12+K6H5AZfOmhYlNPnrdDkmNZQLoyRYkwy+90cbMOJyD5gLisXq
1mwTIGLMscEBk1PTd1TupIse4IrneiIvp0XEfDXKAUpIhO88D/6OLlmpNx/gaqLrhcclnFE2V7ZO
SmombuwcVXtIPGJv7egFhWRgWJdLQgsf4C+Sb6NOVnueLArQO0cBnv5OpuP/qxj8eXqnqeSuNQlV
xGcpGO/ksSYCKVw7LE7toT40TvP5N8dVs66D3T/L1a7j1hQ+jjT6gknIGvw5iNAy2mYMvddMXo6B
H2SxIUxSWy6UcljOxh5xD9pcDN3jZFcipuCEidiTpgRsx5+uXzG2fDKmK8JRTkEDKR2Lhgtt/vz8
ViiYEbYhe0NfbggWcZXPpB/JPXgIgXC86rMPsWACJC1TJXMrFi9TbRp8duOHSirrhvsfLGaRU/JR
qmNg3vrt+ip5IVCZzNvWWFxA5mYxhIt2as/knpeewtnfIwbsQ63448/lMOPtLaAMi99/1Pw1Ph43
nC1uWwzB0QWHLRxf1JUBqdzyXXWRCwrrfc5sWi3VHRD6LViLnKDOUmIDpCAwVSue7pLXs7e0gMHK
fWqBBN+LXv94HG2WwvqaiUcbTyXAbux5hajfOVUIY1UA96OvseODOu+TC9DN5wZVbg1FEQhvAifp
hA9hr0BUb7onC/gtw9EYG6+QIoJ0N2Bc659S11amnu10FNRnSrbizT9fzeOY1f8SSHVys3YzSmRh
vOf0LmNG6c8xX0TOJ1Ice9AW+8a+BWYj1+AMy/xAAvxc7D0f8EH3ZErXP6cwILTsHrlZVb2USEeY
5dvS4Zbv8jCBA/OKBFtXhzFL3EVgEUPN2uH7gwISswtWkia575GOO5H/gBmaDWTqF9EkorLWOpP2
IopY9r4tbC5rVqn2l2aI3ubgkD/MsMb2gFb6pYK2wkZQuwqkU5HthRX7NwHI/xeRgaLmWsF5Qic9
6cRNR0lIWW9R7hgVL1qzM3V5pT4B2776lGB+iXiN3gFNkBffmKFO2S9WqfNqVl43AcX3cqdr18Jw
2ZTD3EqmGirc9fk5DpR7/45lMpPjj2C52VNEXpcloynwqX9f/b6ctbeBZn26Jl4NHJgQh9tyRRcT
ZLkg+eqy676r7dWGQwyMdsR0gFRj3nK6Hh6OWSKACzTwn4z/+pLVpDTqBroxK4os8IuxiciugQlS
a4CqU4pTwUqWiKralvgLWTdkAggelyXTcl7jamanCihBj8b5TRPzf6eCVjD5EO4HNh3xsMjZSSAA
nXWZCI5dhjGlFQG+xqdi6R0m9wFlwz/v2ykhRc5Sq/yauEUuYp2v3tFPpDnmLakzyYrH/N9T67+F
EodBQTa3Sm2eH9vhbTokjgztEVXpMXm/DOgb6J+X2vIK5Xnn+D6hb0jhM+s7h6yAXpWSi9KjmK+O
Xz25PmBKFf4X4ZR41Bk8EAGrsmveskjBfx72IgaLXcqz4//Yb0iVOUQIt3pPWDwtng4hriecws8k
lI5EJTkM1/EJr3B5d4o854AuefKt8l5xlS99jKfcD2BbkacLE7plwytyjMpdUHNYojeNPprPIOnx
RNM1rtOBMffS5uzosO/N3iUYuQ8Q5B1ddc8doM0X9SFdP8Ctq8esM4A/L4teM3G8gZ9TeaOnufXh
N6P1OwLr/AWHXwaDHeV0ppjNfQbgqo3375uqjxd5z5DA0ZcgmaLHSubZq0gXeTsCSrVqgSpXoUX0
byHxN1NNn5T1PRq4idF9v0mL+MwDaRiFRircE6JM68z+tWpgLIAp7qbJlG8b0rhE3oKBS32TX9yk
45lHp8cfXRrO856Jx9+l9iKUb8/Wrn5jiXwpfYOX1t2n4/IxmuYWe/xrFoN9wHDXaG89PeTFp+2p
Dq+SXoP3C0bgSwzJ0vvniXfw6NrUHfmISDgS5lAIt43NwSZO4utVBeWXG+YusAlvlpgodbAxNei6
FKifiXGa36Np1cBTV9Ag4tG5OMaja9RzD05T1ENN2nCiJ+BGzK5HMBEfGAZKQ3/RzWCJeoWug/Ev
iThZZ7KzWnMLAkSzJaQEZf5mC5Jj8Sk8CjR0igzZ1SqfLu/KygwZORAVnQJ27ddFs1KN3YM8+lnK
q4fs/Jgo0eITX8fgYuOeItronHCjrTtmh9szuZXNcgaUiAcSozT+V2zVq7ysMUSmcrV4uqTuFVAP
Rtndq7tZWgcFkvItL+KVO3lfxwt9U/6n8jiennI0QVuzh+RIocg6rFH6+ApWxuJcr2hRX1Ii3PU0
faanYvWj3X7X+HRKYUn2A/GiW5CxxhU9jm/cqBICGhquFAcicRO8l9FC+M6CafwW7+PCUJbAKh9Y
kl+nz3FX2EHs+kI7UBXUmWMKhfh+554slLLV5qSt6H+n6yiAx1VZvIaM/1a3bPfTX8v2uoCb54lV
V19X7blMjeMmLG/XY+4Rt0NDItS7ZL3AofikiaPHqSXhLBOhu2XgW5yr//yMnHzZdJXVhTKPWoPW
TBHymP0eswu9aZiL/KQxr4npeRmBsqLwvvOClzzKVH3CzB4AN1KQIGU2dm54whJfw8VXedKiSlKw
rV88Svhx5+37GMSLpZ23zd277Ajtvhm613buurVOBPhwbTsfdE4LSq8Xb6jPqopSIhU+ykrx50nk
Dzlo/Nspscyibq9xMBK3CuOVccKatSSCHE6ILb3XK6hJiGL2+j+l7wwJ53kAEw+3vMUXxZ/xHXEJ
uvkD2DNX1QYX19VmMjVO2Vfs/7JEVsjvydk6buIVaV+I6d6FxvuEgFjCWMZGyhAHZPigU27jMG9N
HtOOpUD3IzD2RxmzCW3/w9PZbxFIc9uMLlSWFYBKwzBGUHHuzIAEgYYZOzUrqAMjnYMHbIOGUgTj
H4Rpcgyy0RuTm0iR1omeIgCceKA0XdR1oq8hKAyjUx6gZXLABxeLT1avheUD52W2iK4A68YDXeIR
7t0oHAg+Mhfyq3zh5iHyKZ9Rrb9bwaYRP5JknwLXPdPANcolIvrJN10Ic2IXEpSaTMKfTnsA8H/c
O9VoC+QXRiBsWCAVAzRnGJ7/3y7yZthW0eWJ/Am9lwF4amfInGQzAMtDW26ZVegcI4JrN0IP8HcK
DZGIYLzW4/s8GxKMQLDSiNNHey+y0oUSw5Xcxe/4Wc5r3C2rP7IP1c2Z0GU9IoCGd/xc534AsBUy
HR5baMusYmqjCSx4K4+jBtlTtYLPQcCteDuc664apQCHvhYsnZpqR9Q5OktgncG52btWS01Kf3V6
Sal/QZaR8N8WYzO6Iz0Kxo9WxhLVt8XLcI5nqKiOkUv2HLM4g+aoPIycpSuriENS1ApZa8IkH7dv
It3pdiSHOuljc1/wGzL9Ha4sj9NXvRbA293Gd4nU6IzF3G+1oN0OtnqzJbM395L/HJSRpniz3Vpi
ysRfKb1LpLUI9+uj1Gjm0GaLZOoRQMUUjHTP3QRSPH3LpTgDSz6dOsHf5P65Pzh3m/i6Q9tnFMxe
4I3Rc/fwTPc5VqeojEvvXFHV4xr861kzrrCZjsXL2nhFAnPxhBGrY8zRZsS7u3DtEYPvyW4wzAPb
D9tML+si57ehdUfnQs3yVM58X5y9T55ev2RtVJHbEaoL0xoROUUgSnl/keQXDaeOfXCVNZPD0o9A
mETh4JFGyFHniSFspzEt1Xqb3SBbeb1phFkc2bdZSswyuIIuHW82O4WUgliKr0SZbuFwSVp5FMd6
Wj6kLq8HbcaBCTOMfSYveEI2tIKwx9eu50r+XXgSkzHYh3VqZjcLyD5QbB5ZWQ56+ZHpg7aW4zyu
HYSPYkw6lEaReN39hlB99dco600rBcEtP0zv+DBiYZtuc62hpWEM9wwve3m/UrrJyfNW8KouqlZG
Vu+0njk8Pc7QQ7s3GAtklKpA4R0Q6n2AQVVCQR0rfTqeu9I/aN/yx7evJzFQTb/g5FhthIRJvv8p
xdhbTTTnhl+TeabHt8QL3YUyNVN4fhnAdbYLVVm6m2JnwscTE0gaXFSK9gES+w7DzJFiXZs/gBgK
OvL+mPfB36FM2/PjwiXQQw6CpLW3BEmSJ642JBkkxLd/XjKj5+3QYsxEy+rx9Kmq8bMEvpxikEw6
aqPT7OD3oL+agyNHV7dBKIkSZJJPJK35WAM+WYtkj3TE394HRFL4TI1MXtihB7WOeNG352zkUbcY
ASAG3SDXnNDbD8MjxGNCaevhGS7Z8noC7C67EPmrGkns+cz5tbkos8ydy7fGIetAKdrM7cUYRRto
GBE3bH2p1RjoP0FsPsI0TFN4e3GmCtHaKXelEqculcDnaTNcg6FXVjSljO41uviCaCPFPpITajHC
PoIQUsJocPjvf4fMA5DRqKak4vXwpAJIkDhU/dIbpbDxzrqzDEhXc5WJZP0WOBjORZskBG8c913T
+cNjMk9pNUrFtrKH0o7aV7ItJTZEQEZZF2Cgluw9ArNh72/e912UBtFJHJjie1KHsqJlveRuRrom
dCCIreXsh5jdbJ1SC0qK63WuhAEdMo04Eo4hW9pSC8tsmF7moD6IIqRZncqGdMARXlNPwpqpCqyZ
bLnRNUNHckhzXA3um3JrBho/m56CN9XR70Kw0J7Kjf88l0I3cgt3KzZUCYN/IcZ94glTJXVq1vkw
AGyd/CEvt+Mj5rCQ0pWAMtieMu767AGGXtQQzQIdiQpBLIV8ttByMqw49ISOEnbr9MXgVX2NsBiq
xvRjWgFlgih72Qz2xSRRAG62ek9bmxR2lcs620eyeXwx0Vxj/PlGV8uFFV5rIO/RfzMAF2kMNGmN
B+xj/zG418I5ystzAlPL3qu/Ir9z5GQa0S5S/sxN4p2oHjjjmVgJ9y+F1OeaUOhinUmXhcYXgkYA
LPLvF/4p7lVozPR0A+FEIuQ7SJMAzr8/N1sR2ChQW0GwddAPtUrS/oxivsYxSSZ7jggNOaGyDszk
Ac8pqCtG5UZiuGaqLtqgaKdxkB1zKeV0abVTsYkXsSe1gMQDBxgpcqanQg0Tfp4RP40odSky9v6x
fzKRSovDxeipPxXKfADJ6Kuyj5an0TvfQgNqedlTlUpjiaOii825i/s9siCo/dRXy6ZQyX8HTcQ/
XA/yiK8kDaUYyVteRKbzAqvsAv/Y/o7z0LjfRJvwroIxC/MsFqyVRgO0dNJ76Mj5e/8jqc1kZGuU
K+Lb06MZQMkN5PipXPFrSzZZjP/MLKazjoY5UYYFa1QUD6L4PhbHiX2zVlP78av0qV/KQuRM8Er5
tfPC4+6RAgb7GMt6pqepu3ZMfaAiOiRE5YzA206RRtMLpv2H5STVt6JCPoEUxEDVkzG0FVBUOUFl
rVWaGpm0zq39UfCSbv4vnic7pHRiFh9iZ6edCu/8XJ5o8InUFHwlDgf6M8JCzyXiyJa8H8Ly0daD
pMMcZeQSbbeZpsEU7HklA+Wsf7RV4Uuu/QS8RxcO+v9y6o3lkQZ4nM+Kx55r4KLeEhLwqf3qMWQI
exnGcrkvlumWun1dCmRkX1y/Zti7HUHKbCULxlzmXOqe7lDd8DM+asZa8pBZXRRTj7DnTuLXcGyE
DSCYRANw+T5t/rniJddP+5FnBfw/kr7ieSA6qkrCQw2tBLBma4PmwNFO1fAaj8a7B8BQf7a3qGDo
xsjkFgMQLbn5/N/toPfYABbhUh4ilEdRc+Zp2PxEaVWFoyiZsbt3aqeFwBnM8rnu+2quS9e0dj6I
NTd8zCT0lfgLnZeAHAN39w/eOl432F6VxApcwel4gTSfzDX/78/Uk0o1PUCkSM+/nmDn9lXS0bhG
OwtLUBs5srghyi7BeDRSMoQAmf5+8C5b5ZlXqwg1m9ByTeRDpKccUTOXxKz6299UcQ6KtyXXuOTv
MvW12FDZymFLKwyGEhOQvUAyGDZMae4VFrf2i5ACy5GCcfKqImyMT6a8npp7TLtVteYIwFdvD7FY
NR8W3ttrtxNVWqr6H5r/4fSS93Ol2eJl7xOs+fUGU4fO20QSbGwgcay+F6omSLBCTINtN2EA4UfL
QVBfqtQv4z0ur79wE4uqiYVc5cZNzHmRZO0J7g6ug7x8fkjG4J40UaINa0PI8PIpdnHka2V5naH8
mQbhHB70ZmSzaorRTVODqzY5UJmyXvo3hc9A9MD9qg0Ea9t/9tD5G3qEZwIc6B1CbZj1R40TgBkT
hgXO6fe8kTPtgmptK18G+Ne72iOqmIhDTnptQZcDxBgmuSY5K9XUR/rpsXrrQLpD3vfzUB0lbazP
/84uFcT52CVo3BQV0yR2ANav/W4IsC3uUem3QcIp1fZS8/nF13kb3u426nzbbM4ACFRoXOH4V3Ty
bizQ+n4URNVf6hyN8LXTdBsGMsNVNP6aML6iZy5bCaD489Rw3AM14klVm5Qww/I/qKqmbtljGkvL
5aXc6Mhvx7EzRfd2+5GtHeysvk14SOJzeGg4xlKWA3tFIHHvS+nrT9eNERR5pIyEempQToOviLDu
wpXkJM+Cc4PluDkby5omm6PaEz3kVxuS7RkwZYCCjXZsoPv9Qbwul+jGaPITbjR/cFeSfjJL45yJ
BnryBVLk5FIOXlztBLksnL7/20Yx62Q2GI7BGG05xtmhxSf4gqYvnAHJQ+KvrqB8h8WXYR0YJAo7
hFLqpj5vFH+4khpUri3SVeqmhyzSKPpje8nPSsLHyCKAYuVFToCOOcrAKDk+IbUva7T3kzLSfgJh
TPcN+RareYkN5EBTfZvTZ5OqPVmF70+Y03UzaCJt+wv0TrBhz5pxYcxjlC3Hmr9vFAEtjBrkHpFb
ymhQc5CwMtE2TYgvqkR5L7DhGm8uQmvI0qrpdnlAu2Gf3oO2mlOJjlV+M8dytmdGrhVUmOG9qF3t
c0gw2csBjvEXFx8YipMmBhPXd3q/PYXQ7xUSg1lDQ93VcBLrE79gnekIjW65+K8o2TkzRvhmaEtw
nHqJZFWhvc/XptbSKy/0YQ6oSJuPWanTAelSTn0cB/4OhPGjlMXQijxF2DWiGms5BrxPVNb8Zlcn
vrzk0B2WPGZ/a5RSxzkG2O9AGuJd8l2XGJfIUNkrc+2kFVeBHGdPPsgqcPRQhtsY9VIzcdsCY2G5
5HVjJZHLdF/A6qNcnaEF1VhA4/6f+iuMGsC06eDfYIkM4THbc1hJBS5YuKMzxI4LjYn0xvyaXhwI
gznzah90tpyjl6gABxYfbrwoNwMSW/AEaVXy/p+HEZZlrKL0CkG93lpb+6qRLJytU1hGlOG4OyVn
bNpW95iGuHFPez6bOm8eifjzXcYgmmgYuCd50uWwxHahWWF6ygYNG3rws85mWsSZ8CL+G4+LdFAo
G4ScGMhcph/EsXnbM6TgbuuZ/Z5H4JTnbX7dBFjCjib5zkRc2jfvKmXQ+ViPJcY+JlAH7Lf91ASG
2Gup0W9C8PI9SMDnrAsvQdv3Qo30trwZVGrIyJOQl+kTW+zfLpEeWoWDN05PDu39+pGlmTjCwhbd
ELvxEQEmqI53AyhFEgOHxWtw1shZmdjVKKyhC7TqVgIZ1l5hlHP4+IcNszLKYmeeQtJs5+ycpKs1
GMLODu6llYZz9yiWj7msksCqvstWs3p0HYkCIs5puXjvpuY7PhSbC8mdPRELkxrHRb2yJlx7yshA
VbRbLVegQBYo65WrCYP7yhP9RznsSgOvKDDz0TGS/YIPXXh77xX4o/EihTYQ5CBFfbbmY/s5MWOe
1Ia0qVjYTQdKvF1xMJCkiZPe9FHOb3jSpReUHUfIgUo+oQnDC3bflElm4t5Furr4XGxrw82qt4e1
zdJle2QRL5Jls67ZV5oqI/tgfbru9ovTKObVOqEaTu+pPJ4ZJBCWIXWtPRQbKPtefHQHXxxQyIXJ
BGCfFjzwavAe4kji33ADV/63D2hltAzU/6lTZslsTTZcy/JEnUGtmbXAIJ0hrZaj/zQpNBcJ1M8p
/ziEX2D+nmCMHQYGIXk5vBSUQVI4cxZZna2btRE0vSN83riUFxBAEyjldgKdiKcRTavjUyQHlffb
/MxFoFu5uLDPan1SfUvk2wHIqfX/DzDBRq3psfAdqq8i94GqzfCJCTiA5xCOIBILHZJTcq+YnJLs
VSj5wmHIe9R7AuJJADZilKgua9u3+oHYhHExwbLDUbVnxz+w/i99I/Rzc7nVI8C1J9RCNekPBM1u
PZ+pVCgdwcppGYxCl6OxTa//LNDaLrygO0+b4SliamDyQdsuLa4QIMbV8x4ETKMdbw7npB2Rl5PY
WmKyHbuhKXVoRj/LplfqPFASDGNzRFZ9uaUu8xza7nSsjrlwtxBSqAKQblABI+jDNkQZQB/J2sk+
cRd9wlmJE7OMXPr3NxZNymQXix3I/ExbZWb1n7f3lpyc8n0/IVd9zgt08Ro71n/aMp4aNZMsdc/V
ECoNOg/xKDBgQfvh25XiRJ/ciXvL5VBYMAy737g0gylKkNxnnHGvy61AzB6AxyA1G7OCaQty74ke
ohk7zszs1IRaWhb1+I5eE2m/J7fuvhbvVoGBGB/eCKxisIqf/7l05f8v23VGVt1rkgqmezMOd2Cj
Oo2CvfzTR7Hpsch2M6PBgseSVLGgUeYLpiwxkCl4rl28e6SgbBh6Qz0xbRAWBO74RslnBItO89mp
jlAmRY/wiKqmFpwRcBFuJivCQIell/48emorZ1shhFCmmFgLtLWlpZPLlpEqfV76wzFMJv4/SUI2
sos0kKqPxSsw7nYnkIZeXK3XGEMYJP0cdiiwanZjshBgiToKyqOsvd9KTfFOo5j2uyVFfBSBkofW
CnlF+CYIr30u4crSH8i7VmBHPhlYnyg9kwAMlrRqDfoN85Prwm50t41uuG3su0gochZNUFdeq2Qm
hWaJtcFYLPB9WXkY38NDEG0wx4m8VMWSN6tDninyIXgi/giuXa8g7+8KIj2Z1sc8lUwd6AF5FpI7
+m2ouVHDOg0t4T0VdOzeQ4Qv3SMmPuXxrKQg6+dUAn28U3HbaW1tPVoSDDrx6s/wAqYK/IvIiIkC
vONTISJG+/kKS7IEHf860C1z1m+v/YDWPedNfIPWm+ACWvgZBt8ZKWrJ2F88iBPbxMoAIPg5/uEa
oB/E66oHRjGBn4KrllRnNDTgPV4hjwEwODdWRoMM/A19Jf4quTf10SYANbrqevysnIl+biCzpnoB
UBTJu5nhMVMUOP4q8+SJ3kruf+fFmbRGarmE59eL08cQw0HpNIEGsrjHzEegkvBE8nktPWPI6fDe
rx3WjyPZVeJc2fusspJiTtlfO1nTyRT+69PXdUy62ajsz1PhIb0S5jQkFquI/xyp+/e1xE1PAqUv
+6dFTUysDdT2ykJMDzVJfO7Hdp4G9cfDsuFz9654mFIvgrLXQl1hspw0RIiZ+1CpODDkyZ/xbEJf
e3UByRbT8TpSlWCW3FWw2IOJYb/afmh5PYWRsqRkRYmOc8EiUkIa2i4bS/ExKSm2fMdqKrOA+GVz
9J8zlU7TfqQclFtgUXZ2bQo37FWggSHfsuW9hj57DCY/EQGbmcpjIn4ApVfFDaD3OtTq9P0f8Y10
lrTkk6J/aUINrUJqgMuNixLBWYDagQINzgG8wq1ps7L8uMIc4j4HGCfR+yvvMYb77fxRTOOeJbqk
lDQD61AT7A5p9e9SeCyRdZC5gTYOTubThSmRoh081WXdeytLd384EY41HBhdac9hKhZ1KGDSRImt
cjQrj8+pyWS4+J5rI7MOYVy861sBl51mzuprnJvVnUKZI20zGj32CcqNyfVI1sGsXeEigHnQhW5L
+MPOR12HpWJKEI/btUJA7QaSwokPHYYUDwzNxVahWk4I/hsVgs9+jgphK6BVBoj13v6y7IwE/obu
40f/695l9Sr/Um6mShcSL1Ry8D8SsMALVinVaBVEJDyJ3lsXUY3A3Oz18xZk0yortx2hA6RnOmS+
ATs+NJl9N+q9qUczyXAblzzEEfZd+rlfQ+AkdATE6CqkTJrRLmQdXPGxlMU99stvv2x2ruXKfInT
zGaQTYe4dfgz2DkdeNmkj2ufrM3jNysHPlYz/pWa8Vd0/lbksDkh60HjvZLgLauveYtpC9Idwxtl
xFxdHaYCG57aSWyUNxbgl1dgXiAIrKT+hpxn/PCrsr5lRVfzvtLuLcWkXyllsUs9SxpCXwSfX3ir
d7h1bVbzqvW1IBsUdp+4/PkIM/jfaTDMMjWJTx3xqFEtWufhO26rAWoYGRj6jEVxYgfWQISTMBm/
JSU0HywzzuHcRsFqTOskSF6sY4+gd6oBAEQxWPCmjQNHc6EON1huyR0hSKyTDNlbo1aJX1v5qJb8
ROZ8IyaX92teSQEqrTVcX9ploBBIALXdosjjPTos5vDUK/wgZuHf4BUAoZuaIPpLR7ZAnYXcw7sW
cQIA5Zhzw43kfzZZK/bZZokx70UPLtvaVXoy/j5Z9ZqJY7ToRy7PoFPpxcLSUENvs8k49EcZSzoO
sGojbBeoJyiCr1WfDMB9LMJTIcBe6YvOYp2sxfbEL1YhqLzSSlOYeDhKM8OoD0kM/L4C1ptOOIzV
X81P0CSw1CtUQ9t1MRlggFGj9Wwn+7MkYZ6OJ1AD30Ur0Hl4kNoCXk7DT25spuu2E0/KSUts8wlk
XGhV6mmE8AQEBpK0I58pv+tInaLfcH4dbr5OXhhEpPptSrLL/71PdYAEGqOlszf2MI2ggDOPi/5r
sxQdhKUaMmb4cIH6xQF08FegZ8IaE7FdSJlbmqPEC1MXNRkESrLyKy7ba+vs4N6O9Yvll5PkmtaR
RcjnO2x5vjtHGGfRbMHTK0JldG28j/TgJqkBGoczVr7O6QjLUANaR+/VrEvKWAY2cHjrsU2z2sRu
6/OLSNO+DdNuBdfTefNpbEU05Npza+GVcKBgwh1AmDC3hx0vV8GtItRcL3g+T7g1clJ4GjnMXnuA
alQMgCQIPlD1yeJfRm/799ilND+yo9u1nX4rCyykc4jxF04W8erz4q+8NCSEM7TZnTZ2cH96dogt
Bu3/6fKKn2qR04C/bh12gvKprxZta/oe+It/UTwHWKt21rxdaBfRG3ke/sWUiBUwQei+9+ANV/7+
iDoKok7HQYtwK0aT/6fsAjvwEQsUUweOG7nhN6Zq1TpDjNmogTooX4IjTnxD6aLWuHguMyB1Lsl/
zeJ3TN8FChcl2GhNlPuFIYocoxwVgkEFlQhBqbfWpixVPVRWKrGITWNCgkVuHFNuIopuefEXdOeE
05iceyRCA08mrYhfQlSkbuVM+6D5BdKKqendH35Lppl36yUn1X2Tqdtjr6UNz4B8KRUHo/Yrrfby
zCpWckvfXGmYhFtSNW/SqmpsY7Pxxs1CBp6LEKG+GamxQket7U/pZTPE4zNAxo7gLZ5d5sHGub2n
4VJMj4CkujMcIyLOlZFfgNFgSKjLWApsOJRrsBidTRVZsxZdtDGIkKxUnyV9qVnRChccBamNTcq/
MRUcTzn6irzd3HWyzi297bhvGox5j9n4ZNE0jc3eLoywSrYlaLlojRwf2ucyUrEYBho058rGN6kA
HsNjjwlWJ9OZrJ5F4IGMxDw8rUex+FO6nKaoDDEyyHhqQuH85KdMFU+Yq8/XRBzJ3zStG/NyfTzt
bdxzc87rEn9QOsp2zivwHmEZTLrHDkCuMzESTFmiHAZsIhjV5DiqVAGaYppvN96f/OuJlOGrCJfn
IGvtpMG+emMauWzGOKhZSOwL6ZFflherH4Qmsb/xiAk4o2CvA7wbrP2FmYdxgtAhOYUYs74XrBrP
QD1/OYWuB8t1Z7Fhk3We+bxn5yJJbk5HOSBmOxSzHgY65z4EMZXDWZ40YQCS5Y0h1ZCDryklSgU/
iQhpKFjaEvxOZZyOhyF1UORHXZw65/Lzg7EAA5FeR2kl6igQsgRxnrTWE9Uw69DJp902zCo/xovd
SAalqsf4l4zrGAaeifd26QhXQGm8+XfmvNkqpqDt47dpIKaX8flh5ZLkBqiC6WZSYxWJeXq7wsrQ
GpEXxAI7YDspXBm06wHx7FeYZdbPVopQq7dMn0G0ZK0KzS+v6Us7OFPds4OAB2OQhWfQRsQcR+eD
03PQ2jzQHQ1y3flsfYDybe/d/QAiHniI1yPpWdw3gRMhWSP1Ed+qHtAYYMIe2zPJLVdeKFfqfo4N
Zyq9bhWy8j3dqKXzBgLdw/rhfJ8nJM2kmSXsAmD1+2PnOpRadAukOXDZYrxzNBFgyKHfxqgM5ml1
IrVbbdTTJIKMyv5ApIY3AzUmlG/KdXF/V5beJZhvoWOXwCnJ+8ofKlXtEqjJt8OY5SCrVRRNAXd3
zFzWThAG0mwJk2D/UbYRFwNP3L6e7xF9ofjW51shIwgNfecayd+TQv84NerfTt7mpWvSKIbU3igA
ltV8BBaCIqo485UslD6T2oD2p0T5rzWnlaCK9WDUSe27BcGBnc+Rgo3he6ysQEHLxD56yPSWFwzH
rNLja9uXMQ3fak9YsyMivUWQGAaaxYGWzWY2j3um5I0B9I3PRHHUlJrs+ItcxH4491cdyMhQ8pWN
McP6WPwqK+Qj3oU9k5TdFNz/8emoIQcEOsDARxWDhyp0x4eLiGWjTlZZTTC1QDmJ/rH4FgUlkLjS
kHtddxSBe78wFyWPXJQFNho9yHLNS5gIpi9C0yWL63VxbNLOkkOKioDPG8ssXGsm9neEAU7Ouvg1
c07IcC1NusBh+kqjUZCBWywGHD43/Zcvjp2mcqavSCDYKfZ2EXHa7qd+yDBQgXaP+jdRynLG90DE
0X0cxP/Xlby0UYsWhbcOE0bYp4joBLQsaNKmZpXM0wzyW18jlfLWwp1UoZzeuNtMN6sZB1r0RGrP
vFhHUr/hm8aNmTQ+7e31QI4KjuGXcOX4YFJs/vtYxDD1wNtneUwmgL4KTRmO6Ccn5JWtUo5eOXri
G0Ato3oIQ6qHeraxv2uunbKBV2itMuMPRZP+35FUWVtTqJL5sqVC6pGxZycntLJ+Z+xYmVhTwIx9
KoBBgM1RQKXELeA3gqXBJLe8uikgcdWIbI7uvf8gAX/rlracaHCFNi8hN8p2f2KHMbmECNhkyf2/
6l/fiPkVI2P2ATP0lNbIin9dPEIxXHtwC12VlTnOZPbswtfuQCCrjcshx5rhDdALh+iibtC8cCcH
ROe1RUH2RGK9gkghnKhCx6LDJnbizkYl+sP+W4dYWhR/6UwqKhIroTqsaF7E/kuQW7p6ECzBE8Sf
Jm1ovPRAqwvsFqCN1poJiI+g5VXNcgENb9ILQywBQ16J3qSWiJGxjHEpV6YD2JDUKloH4B3LB8Ar
UcbweKPdwIkek/htVoG96Y0EefLLvDnotg03BKszr8lbbJCynAnKKmuHa1yyQ7VNCWvl+fs3sd3/
tpPA6baLMIIfrw19KvMKqbUeT5rGyDyF6lyBg7uIV8bYVIC/plT00ByzrNzbJgReLSDarhpPZTmO
m1un3iwcx87CufksfjFq2A/QJOOAnGZC+bytaBPSGNJzuF313b31YWKOuH5t8FulqBkRDjtaUqzz
Czok38cnnx2ip3L9m4vFcc4YprZH86qZ3trU/RfIdxUvAAcP+qzGmAOrLdcCRBVMAnNw4csouwHW
hzsHaM9VJUWBvO+Z2ks1vSxWxb0Pq/X5GiB2FFvmY8XEmD5XH9qVMsquHlgs/buX4aCZI2aMRN4K
sB02Qwc0N2zAMWJBAyLia+dvkNXy43fVDrxDetUCaJ3XENr7t1pu9ArkwJcnD2K8zck/DcC2Kv1a
m0lviniJdp9nfv3wKGrCjtdChuLlJHbQu84GzhltgAy+bXONqV5LgtjFBeBITzp93fxu1vPDYi7t
lzKsGZezevV2XDaY7ulr35/7GQSluxmGTk9H2t0TZKaFK/n+qeBNtErdZpP92KSHJ7lQVL6VQUGc
Bb0a9xRsbnrvF5oSKiezV+Efj8x6wRcueD6AHC7HZ2Ao6SeX9VgKxlCnU4oAkDxTBNGd3HLCZhlX
w/xGkOUDE/mZlCCE3rFjetxlmu8uY2SzoEEI7+b4y7dnrKkEkhYaNxq7rBVgp0srWYMEQ4A/ZWZ8
geAQf5JRLJ3K4JS4frhAO2lqVQqnwrmef9ubkPrAmLlGaBkwaaJZGBCCvepdL9J1Xm3w3ICi1wUG
be0+zlyQ/SoAkXWMpgL/5bNfy/yHyeoRpV3x+TX01bMGcW+pzmq3mG4A4jUYN+kTTRxI77WRoXUL
yIgRPlvDSMdk9Xxdq6cfugX6ASh/sKDVh5+medsj7neli2ip6rHkWxeAI0GEw5IMoXr8VMcmsBET
Bg5SZ/g3ROTYBBmGDW1jZ6y+4EQO1MFxrcT9r43bS3ZdXPMwmGzXyvGUlKyE+j/aUIu1gXPOBGUh
6ZRr+Eo5ZE2vbMHrpg5rbnxpLpZC7H3Rnbjh7QDk3GpAgEkpAgSCtek/R2qgEoRZu7+4/0B46T9z
oB0UTsByBOxZdnhHJTruL4Rpv3e3qmUEXShdIEYW3z7zMrTkICu5zPXrWfo/BPJ+MoFHj2G2DVSK
xF9c6WuN7rJB9Ec+zTWzEkipHsD7xY1NuSeIRunZNCu9RfoQ7XNve9MrAhSs6dtmZlw1IijokjmZ
f3XJzHwDvltRMaYedI6Kf2vden5l8Tq/O27BAk+3lCMHazWjx8xgo11pKKwCH8s6bwF9L7OacZod
92ieTR8YH/VJ/RtzEtkRlu84rtV2jRRRFL5XZSbQAXO1YOgwl1ZVxwNnZY5vP8r9Hn8oR/PQuUwI
7SkUlYtE157Ref9XFcB94ZnmGRZvgjMnOe7WbDmd8IX1Tj/n44Ui0FidiRvv/4HrIL1ZOEEIg7V6
dTuwuUqKNVpZW7JmcnSgSS8HVeHyIRaUWTH6sZvpmgBeLgMDSAFUxX7XDl1QRDjaBBrzSob8vF/M
ZWB/BBPugM489evzK7pZYYX+RKqPa5d28xgrxyr3z7YJESiq4EMZlypTGTDCLR5s3YuS6nRItq5E
021RTmtvEuJZv8d5krN1wAhLreQ4FdE6ygxFWErTWeVBfKy3Bk/hEqpQ+rYJr8pqLwWAcwnlVJDQ
TGiAWhW7ygWVVAU1Ek8vCfS/skqWK/3MByFHjCg2vy3z17OW3PuQJ2nciR5e/lc4YlSZBRCeCHy2
SfwPQHjmYtuwG7HLjjfnVzNYE9dQi5HGrDi5rkqDaK/dU/qg9vLiqvUrpEjbxuEd4LnZsJI7seS3
OXUNqYaxXZCBYX8BfdlbovC0lsNxFYiRIlI4ugubpNWVr57bCNPviH7Q0ShMDEqeKt6tEMFrgG6q
zo4MGfY5cDJXCSnV+b9aOJLOsxHActWaUn1KrYCX/DZJ2GQiiNYLRJ0ub+0SvSM05fpJtbrJTNmt
5jrTzp2mvvt7RlxSw01xbW+QUik10Cw3pqgxiHuzWtI00bY8LqCB55+4DquTBPhya21THSlKKlD1
VhbbpaNbQfFfpwdC9uifOmh4SqWn8eOUbiiqTcAABT5VktfuS3AIHDlJBHBrOagHJKGbw/GyUm6G
O0UAoSIm+vl+fhhr69ZGJyjqfp/R8lgu49oVNwtREcTy73jy5mx39VwLE4Y6KBLdfCdDCPvprZAW
QCI1vwxIxDI5T9WPWU4fF+mZ48o9U6Ilo4XLwngG8XcciUv0Lhaz5rB15Q6DKOg+LFrQT/BetEaH
ErnUVYuF/wKyYEqHnXDYZUUvym0U1ht2EA5kDejbBXynD7HrMzNwnPmNDMNj2sfZQSI/g+Lt9xMg
Ye+wP8mLooazMqg5jkcNlfFOzmyOPXfV3eRvr2orl4PykLMPEoB/mVlY9BqN1TfzJ2E8mu2rR2fd
z0IUKgaW9pBxsGp+0yEp+EL1Q413fRQDtlpJPiwNipQugCsDyaXgFOTCTF/N2FfaptiUfiWbqQpf
Qc+hnkaZhh4tvGwRIldxvHHUIGJdNyIjvHVasIpn31kgH8ytVhmlsLtPh5f2i09E1+E6DNqgh/UV
uK+0e9QkwJTyD1gfcE7mGNon5r6V7ElkS9W2ZudaBHCwHwPcbd1U6K4RBGhmrX1+i02wPmDG5kbj
76te6pumy2PXi5xxyK/4FsOjq5Pp13udOexgPIv7mrVPqYequfBjBPakggdskzQqGNaUzHQHJ7po
hR7l0U2WuyXdrHWVC4loOsUtPyL4RvxfPacXciTmfdQOXhZsq7xMO4jb32AGaEdAqiDHPI6pE/Xx
km4RPzshDycuvpLAT6ULgtjJfXgxTUqYHxIlhA4wcHOVTXkkniVw9VPtzPRg61LmpsiHj8gnTGAu
KL05RilO4Zkq+lbBdUoa+sPJ3Zh59PfOJUpJuPLxf+WmmExwJT7JXoEGrNqLyzZ9XyYMEGZFMeA5
jCimxRBhrB16jkqKa3jbMzot1BPLrGXfOVALoQoWahB24HzEjs/H4Q2Wy8ECrdAu6PNRNiVIXDkD
e/59KFpKPHjsAeOxyUfvA7tfzUtfeO+n675N3sUxOFjw+w+ykIgmNcFDmfrk0o8FrRlXYsuQTC8o
3Lh01PbOtyitvw7GRkG/Cj8BiSCAE4PUlPyD0ZuRywvqL9LZOLxDuS6Gb9LMfmZkedVO2jxT5Q0I
0N+jVcdAMqPsoDGR4RQRkMmdP2JLPQ==
`protect end_protected
