-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
DJk/swuCDVyT7+f8b0JoU2Wf2AMngvh+k/1AYiZNeq28bADofj1HxTqZ2Fv99RytR6GpLOc9SZuh
oTGHKLnkwGDbs27b5keOc3Ap+U5dw9HWlRt1+rDlKJrxXdRIJE7Oat+vD4gAqnh++941Z+7jiCZF
qRL+f/pUtiDccipuDh2P7xjOVvuQDxe0PObWNKvNcR61LeU68wsCjHJYyjYi70F8mdG3eSEKb0Zk
Agl1Wmq+0jTmIkXONAIcgqsdjotEmGo4lwGYucFfb8FilVPkszmDy8aQvqmPO44yehsumgZAh14n
gZyqbJADzx2TR2Hv8N+9S07BJfT9WVct455cqQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11888)
`protect data_block
eGr2w/25/viiWvkYHt+DLiwR9tL6uSsI6cmsgEM6fh5HBn2oY5o44SjEZwSCVaznXzFP53sp+0om
kwcPGfWwMT4BcGzQ884Fk4V+Lc+4oBTTEsAY0ZG6qRK+85WVg4HoHh+t+/C9VvIQ1ZwvdS5Ox9a5
nyWeUe/0gwWyi7aueMAb3omQLrBUXiuoXczHUdTQtO6wNvBryxtvI8Hitta3dokUdy9dcGnk/+Ce
xewivDqOfkAa/DQbqRAgrARCBGZ30oQwG6OZFfoF12tvOmdG9YMLrGV1dp9nEDx5iDOht4hQ6+5s
CjVqMk9jFtbbjiZIwreKCRWVYg7P0qN26P9W2Cy/zq4ZxblhECKgVJ79p4kgI2TGQNZuAJxCoZ90
LJwY13GzQV7IUAJQ0vRWJvAdc8goymR1hZfHQ9zVjF3otvoj1VWZYx3I+PimKWnSfORd2UhG8IJ1
oCrRqiWaS/7y+Rh2yW+wB6r6/Z6uCsxDFMN0fcQBhNZDjSlRltr8dSH8AjzARnlRLwIsZBOkSW9g
8CAY9JvLZJzwDlcBa2vJ7IZTVZCoftFMrPx0kbwS5ANrLXjtiX56+09RNh6/V56yxo2f/h46Gldm
lrzT/UIsfv2mYK5Mwsc0+vKs3bcrMszLzdgKewbSEOu3lsO8s0CPiwR6IYfldzw3bhp92lFtHCCy
NT77TKdnbacrzZ5vhm8cNBeIJ7/mpV4A6Ovx1FiNAIMYz9VCPO/9ld8ybU82u59T8u1Msl+XWBK/
TyBeRVgKxI4wGFv9UrGqRcSMrv9md+1eAx++PfkPzzlLzK0HOqtJZMSjLWKieAV7g3hOiKUfj/JQ
81gzO+sCZzbqC3aIhfSCIjujAq9h06aY2yRbP5qtevSwOe0ZCi9Voi48Ni4I6GntOjFXHoECiFDL
TnvsI+gzN6aAE4etPOHPzq557r4kayoAi9glW0J/TIwzqPOudJ2ETPB9MocASm0pDL4UgzWFev2g
ExeWaD8JG+hlQVpbuCCeCA3U86gFSG4S3F78ILqf915TKAeOWM9fNLvUJ5dMOnyqMR3vKVYqDcJt
eiCVrkxn+7Y1wfYzShtdkXG7BBb9f9au9px5+IpeNFIandk+Gglh5JfTwFYJufDaXModUsv8GA4P
I8G49ZRZXge7mgDrD+JrTSGQZrF4F4uIpnqxUTHjtD9reLBNPM8qTGu0nsFSvTa4V5geLjwJzL5t
N6oVzksxRqAYhcZi58wATZPMbRAmBmCxKvxFiy1Hx/r2X/OZbflBkC2zd1NNqgUOR951m/YDU05S
0FqPbTl3HzDLldr3rDlWhImSZuu+uqxJTqKqlz/TK1hM0AezeezdGvPUBcSP0p5367qSYBAdZKvf
SrWp7uZkiIqxQ2XXXUXEPGH+db6VlJjxaOt0k7FYPxvMoUB25Mcd6l/hxNhe9FCsTWbaD9G/yTVz
MMCIO3eIrHJaYJ5shs9ofL/RBiUMAX8AhRxVxPA+TZMCKZ6RkWklYnUitChbqdtHdIwkPAnBkn2x
LMPZkjOrXb8fPqaExRgeP/S1Dkk9MIn+f8DLuI5TczNrh5M2GLYyRmJjl0gru6jwjo4Uc612Du8q
2b8m+8MMnUqvuIzzR8n5urty9dkW+h9idiU7b44iR6Z4jj+zz/jzsj1xrKmSwOx3X7/x5JStwT+1
ieKrr5q/eRU/n2XPHcUbTbtpArbSBZSQe3+xd7uuct2OVds+swqzJi+9m0RHNizqrj8zs5gSAJ+J
CR4ZzpuAyzAWees/EAiUHhqOJs6X4jgqZcs++M5/WfXAR6PqKMrOGQvfPK07J63iiq+uiCWJ2IxA
bkmYDaZI848kQhKQJwC18oysmvcBsLmo28tVIbbXx3gOtH7i3MMM9IUAM0DeEM57nhtQOnmuykB+
HR9b2cqJX/8D8vJeVqLARO1Vi7/IfYemTTuTte50FSrrk/tCx+QjsAf/Uh+CeaSUC34/sOmzwXvr
i2oZoobCHxXVZuMLyiFNtF78tycIVGgfqobD8gt40osqZ7zUoCxgL/w/mNgvZgzTYqIbXV6kyxZn
1rhErmF9ifSKIB0I0n2LsnUeO9fBHBI94SoAoQ/5XqGBiYe9QZPse1hImBHca5mmoADm152hf/8u
19dwDAEDvkUjMyNX7siGwBc4qYSrJZFv7yc6UX2b/TuTGIbJAWcDP2THiVFarkmF1YvwwHsmVXMK
zfOdhHZYdbg65wnOqtGxeZYzvhB04TFgAs0FvjSuEZLzhHhd1oV4nKjyvVcdE3tJr2jwkiw0CuLZ
LBolsomDQI0fF+RksGOPMEE33Iv2xOr6xvclGeH02d6p3yN6o0nDzUeE9QuKtMbOz4bsZKdDw+IO
/5A2iEwzjsg4vf7P6cNIP+4dGbBs1Ab+YI3ExBlrG9gg+mgCrtK390Olafl/RocZkWvt0hwo/Snu
AQwvLDHshQPrYhoUHqdIAqN1Rvq5tBy9P6XsvMqhzWGnzONe4y/ugnAFLMr4tnO+3nvte/8LUZMl
xNlmcP2RQnOu1cv+4iAZDeukjBQFWrJhN/QTqtlDkHBNOKMMn3eDunkrAUV6moIOEfbXGd/kKYwn
AiZseahya+RlefjG2S/cDad7vPF2Kv9q+rzk3NP0aGkiEx7HRGWgmW0DJGTfPChc63IIIqyd+QKP
cHSOPApW4r/mef4lWW9iUpuMBpp0NWft+2uFsI39UBeoHvaofuCpgtZvn8ad9pZ5CdTCgPkyS/Zt
N236RnofTNBWdTzL9VOC/ruM+rlM0S9M/TDvq6Zxapo5JePHb/h3+o/UzYUeBDT2XBpGQ1DpfMgv
WUXXeWNypYpVnoXFWEAORwHXHgwU9HnjQlxa60m7VwSxwWAVyI8rXHn+hhD77cSZMM+q9mJAWJ8M
xKDjAzlC0YU2TkcN3dGbjjrZXop11CFE9FHEDbBw6sWXp9lDmzT1R8l7y9f2g11JWOg/2FdIDx2B
OP56gxyjb0Q1kthsYBzyqTMxTUcpEaI+OJOlGX+tsYhzx++Pby3ZJK1tq3uChemusXe8kdWL797x
SPTPcS7VJqJWeiagv+H/KqFJiFU+fZSSR9EO2wncbD0dmj3b9n11pm+RfKsraw3F4XMm7PwV+ngl
QaHPThGSqfW6kZAyNHgU/Vyu1JyobrtqIqjZDZKrRnAtPJDkSBHR4k7rhsKHRJ0g4vmyktVtIPQU
bKWFGqSeb+rDApan/YAqSFResLqVQn9leiMXFCXt3/iYu6NTl0pfxbZLUKLhY2AGCu5ttFbyB4yV
9IyJFXHSPA4pxmunon8YCtHUI5p/+8oYrzcTGWfNkvMSdn+ogXymsiM7q3axuRNAHB06iL3xSSwZ
rsIWpGitTN/HpPNKimwX4oEjW8Ait4raT94jsxrbq2dkyNG4zd23aOTUNOWD1lZgnVKoSB70bso6
XgHri6XIw9dfD4Ob8GHxs65mWS7Hl5NLzbwq5Sr/4dZq5pGafCHlSL4MbGJCfcKacg1GG2zyvKaw
pOroh8lxP21EvHFNdSpeHYASVdx4z8zWYMWD99C00zH31gzbVP3F6q9p6BVlvn+kGaUlO/aJ7S2r
YkwwduF/GhnliXGWSZyq7Vle38/4DTzJo8MBytlvQZ1wF4BXBOyJ4pUjXbUYjPWi0/mMIlobI2n+
HFUzHI+2xSzUusScN3NAdejEfUt//yQTT+Rn1w57dR1Itd5zB4YY6XCWJGmnqJDrn4U/h4sltouQ
77334Uom2+bz7EtL4S7zLvvVTu4okpu5Rabus+tff7v2VsrULANOYlD6gt4F0zbwLDUvwhT1lcFY
ICBIQXbm1U45IkI/L9KwCgW0o82cmCoteVXw2WRi3hGFmksUxdpqKcX5Z3S+SsM4b5/S871WH9Kt
r3ds8Yk6ohbN84EvsRKGjKeuNSjLyvcu/60ntb04Bi/7wPCnc4eA3Z0xmvCY5gutA2G77WLceYjW
aPkF7lTR4HJ36HyMZaYpz+/vxCkUfC9dkrHPmvuMhPollVBjAg5UBmDSl6ku/GhDaDUC4IGOOWDk
+8XHs6z5/k1S1jR72I3iBv/Azrs5lcPTWRLofPxwGqxMfciWZ2RDSTobJWpE7x/aokjzBst2iW70
VIwzLCZBjBzdXnpa+h8GhXAp0XJ+tGuEez7K4LYagMUP9YQfAPyYbPWdnX6Im1RcJtRWHJsOC/HM
ymQh/9kk6g/rqyxD0NVFMVpWXMAj+IUj7b6a7qYEHEg2vsOKlw1+THrApUJVqBIetP737zRZL91O
Udgns6T03YWyPlkR8/OAcejzT/wb4FOVYFHFYX/I7kUBOaR//jtJesqK85VVeMfvJFHFSJP1w7L8
UIOusk2OpDp5kr6qDV9+9ofUwXmv5T/tzb4+8gHZgm2bLoVMx0YBL9GVPxKpcC5/KHxj3zC7dRpJ
+EIvHtJDRRn7sKlStrN+v1KtbpaO6vrX+hXhrt2EqcNXTkGKBNkNT1tOF/UPGW0qqr3BIsE6Rme8
H8oDtO52XWfFURly3hf6PGe8VRgM1iDp/3FKve8Cs0aaMG/+bV3JXGrFFooKBXoNqvdR+v54tDDx
12oi08ePbPWtli+vl/iGyQ/L9R7ewXEsTx8ij06w168F9e9g/SAOenDXefIu2qzYcI7j/vR6Gbd0
8uldsF9fwIL25A1GRyRRTuh0nphOFlovb7XBQB46aiJ3GkOAYXWR3lCK1p/x9neny25GuUEfsiF1
SDiaF8sdSnVsX5o5eV6vLYw4Aw6JCBUax+yNdTnMKaDrCsy5b/O4TQN3A7a2jlE7X/p9ux8wYfOi
isGXhNoV/WXqMqVMmKkk+2cq5kmSUyeP7qfeDmJh06QmUf3UJmR4yHI9PfXKIKJ3hfkRfQzS+Kwa
zh7+tTn9awGzfCy7lVh5R/6JOcg8WAMZghTIusVBZSSKIicMIe85hhuYVl3f1gisU1pzDaACzZuy
NMr7Sn3q+Up7Xz42WRGyl8ciXTCC5oBQwWrUffKqZoaTOGvS5G85cginyEPz0G4vSuf2fNVMvxw4
OCOXWIL19Q/3oRb+pWKKDgjLQ855Ufm+JKoiykV0yDar0Rfhf6yJ18k7FTx0w3CTB9PLYhgUh529
jcnUslEwErm5kd5SZlHq77oEIvKYxGyCBHlL5ieuYRnNjbSvWM93d5ScZdYrItnARxQBCKp6ehTp
67aYhY0pIyFP1Epe4ZQCz1fvNf2IrQOHbwplnO0u/sb7+cCZwEQD/ZCPuMFyoD7Z678vci0LttFS
CtnsGv4trt75ODtVqikT1UL1maKS3WbQQnp9TQD8PLqM8mu+c9MdCaax+Jbi98exyZqc4Fw7OVwi
Qtv80lL2yzP9BVvi5AAw02SWGaF/vI149muxLhWxL7s/Q3ycKlg2XuxbKCnS73UF5B57EaASw7Zs
jSJYEaHm/wYYtcZe/KFWQZzLKrE4p5RaVIAMMLf1WFuiJZlRmorPL/4mxzr2cKOVjb/bmUdGJ9qI
UWjAhtmdN+qQ+qnPppmYTQWl9FWgCXiYtIuRXKiTs+XmOS0NbwwwehH1gUbFXdQ+Bd7s5KDt12Zg
awXotyF1cjdPHJL1h7Pyu/uIteZTvWLQgM9RfeKePH7kmrN/4ic3cDOl5Znfy6DbNB/d7H1ktFx5
CHeevEkyjX7PNmnwcMw/xohWc1hKhVbxp6w5/n3jPPSbDYCn5FUpVg3dpxW2zeyEGz4I0nI6rD+6
aZi3xgSgltX4BUkxrWbo5CQGBbVkgf23RzPiJsFEdfZ/4xWysQFZcRd9erugfUFPOSWh/X9gsp6R
fRVPbDZjCAUD0zd1GI7TqpjaGwKzok2FlnOJh6FLM919ycnCFNb08Mlns3ocY5kL8/Io6v4a/uL4
XwxDC5zyx4/THRxxdncUQkvgdt4tezz4ZjUdhH6V41L+saxSgelnTyvyox3HTmK6l060JqquYy5+
gge0BERST7IGJzIfJb1WhKS+xDSpb/HgHQJxGkH6TCrNUSWaitw5e8dVQUo91ulP9dy9hfGxP2Qp
Bev2G8OXnS2WAqE+Dbs07Gp8s7WJDfdpLY8WbN7X7rV6cP1ITASoQRWK4Vu4bxWz2E91kQjbADD+
edoKKNCWUTh/vcxhtTzRcstr2NBK/p4kivDdIgASE5A//7qXxzmXdRG6dPmbVg9p0Z+jcNSfSfuV
WyJKbGbyhu6N2UXD2E73W2o3M76Oy1oJ5TY11eET4BKXbFzx8e1Zcqz/iz1TgbP2Hex5Jv5vHS71
khfEXWe73Zi01TULSz2OhDYK7wEIEf7zOTvRSn4G5rGfQ56ISwhTStLFKgBPYueNWROIDd4/ZGVX
+cla7pPw3c7et5oUjp8XYoPVDiCToo1XKhx2nCIC0Emr+jcjYE7EgTSaP+9IXRdCSbPPLSNTemsx
9qjOPTIE7v+rDXo50XKaLnBDYoV9BcknmoTGi6IGEVFX3XW7/txFCsJvtZ4mQDQ5KJYBdhw1Lp4d
fTIZcgmA51SnzVQ6+VNNZJZ+EaBYSMxNfmpgL5LvbWZGTFURqwh2/BiAR0JuVbF8Q6Pgzo99fYTE
2fX7Zu+aWaRIhnHVMHDiwVbELigHBCyedU5GbZewCsE/qJF73q+SlG2IlBBUnSiAppO8GCBaRysl
NYmxr1Z2a7REoVMDn7HljJSExXa4TXOaaF2YTVGbHqOSOORQaLJFX8kwdXxzOCxO988EcyhCZfnQ
ElNYt9AdrHTc9Mi4rAtzolQaYr7kgRLyPZXTgKjfyOKN2cqiO+n5F4d7cNmu/P2e0kfav3Rd45Pr
p4kW6lnwhoDLiT7bDESAJwbWbx7/L1PAxPw3TLUtcSEqvTXRN79EzOgwpGbZxyM0bjeh65G0Zhy6
wsk/8NmfTPxXLwpG+OsoruvFSsjJx51n7Y3HgcYgVcfM4LVatHlGvAHU/CG1jBZv/SlLb5CjCQVq
RaSe/rEe4MOcKeTUwl2UJxu5taGLcuNldRODSkeKUcMYX/96T7L3bV4rQ/FnOJJ9+cljfqIFy5Fw
bAkQ30asn0E/QABySXmQt7orJtEXmzJiMbVffBo8TEs4s1PIDPURdvDzj8AaH8wdDRbgvqu3p0wv
9Xyh76u4Z6QGrWOZqGtwOK6kk4MwhKi19+WF0yWoyjYBT92Yw3gDv7EntQPnSoun8asV637Nrza2
FK3hWYrYMwmnECgExTNX90631xLTi35xUIngR+NRPyjvzfOBtrXRQLcr+1zjyf/c0e2zdsKjxHEN
fT3NmRpLXS0CiLSE/sbKMxSzkc6kVo1uEcCxVEUPryiFTOTFbZ+mXhHKYoqy1aNxVQmYkPaKfSDk
DSdTXF/zlBxQs3noZSWyUq9cTT1YEqFNDIUsDtB2T3wMXkpzDe2dlksOh+vSF2E0o002MS8tucno
RY4VmpFCa5o4qKCxPO6jlEjydWqsh0TXV9RKcfUgHyrV+fknWPbPEVOG5oE57Tl0VmPkZUtnVSCg
ZdCqbCysOJKIMPU+KX9kq4aY6yELsdeJ0U1F9wOd2fc0zwv/GoVybO2GElZMZVcjcGIp09UO5vIg
6D38FPy6LyvuaGPRBYIqs1vBWsy+m9VdzbxQ23Xb0sXN2CRI9stiJkY9odzysv252mCHWIJGxbwa
KC3jOBfl/9k7+UaUh69AGm8ikD3oHI4pSlAZTLgklYTL4DOJH4b2yNCvH6omPsUMWgMGanPBv8rZ
0liC1dOBNOwTFYiHrJl9kBcVWR5CUN2W3YoPSF1xneeU0Z/SRpZHXVgnD9RrH59SmFCzMcyZdTht
mKdb1ll5ycQZRklMm4jKVU+He5/9Gi2Q9begooxgcw+JZ2f2s+cfHyXkzhmVIu88gfIrzu7ODzaa
5DMzZxpbI1sYnTVSJKn70fXtnQ1cGNRpynAPnBRD+4OMY6ioWr4Em+HqyPZHzAqzESNL84T8MLRA
buVs2oLM6NwJYWqVqses2uzM19mDujFwrX6IMCEuz+hu/CpfZ20c6NC71+NeAPdZ2mmWXAB8glvF
xA8FerpvRHJxBjrhPhJF1lcqAcjVXpVpCBipFjNuNnKZPNYH2umeLXNiOqTARyxX0cXzBL1JxbqU
JgvqClCVKHHyw0/6473sLXZTKwvmxgdmKV6ejnBu9r6qjIU8p7cd+1ptc1JmmWXNWBZLf9qad8Co
R72lWVDFTp2vhvkx3DPBxFRHogDZvAaBqUIpmkS3GULIrxADbZ6Qgu4Ybb9/er/c7KXYUgablsDd
NJnoOkWdzdqDWS2cXoQZkFoXMeSu5sqAKtreQC13Oqi6GUBpowGMg5fX6HT/YzCM3aTldUY9m3Rf
tiQ3pDIzjvoqazFjQHgdUNxwbbj5b8UtVVMb3OYlWQ+OcsLQsXnmLKzTbMC7jcXyvn4B4gyg26Uf
3ipx0xjwVgrntNs+xiCOH8ICFnDfwLym1k43bfrHBVXIMElewX0SNCZ2NlQ0q8fGjYNdbC2taGAK
wRtFJw/xKmL1qi48mpzQYJtWWCxIue38N7CUqAHxxrUt7vkzEoJkqlVgkU30Q7J+f4ZPMKm85Kgw
mSgwXMsZBs7FOcuDFATQkkUDi7qYO1uuVKqft4o/0cykVM5Ig5iUE+lFqlI/78YcAGZvAgXJwr2I
BLirQlVYDykJJ39bwkq2OEWWeEfTjcSBy4olvRGALTvxJEG9fLx6dAoUK2QUEmte7YrIooo/AjUO
wTQPDQO3AFBuAhKFmBDRIKbH9mVrlLs/0ykVvXbRAgRFPsogS1ShItEeU5x2PjNmQ0bZKxWam+N4
Rl5Zuumr/EBlSxKkAnOcUNrkQrcD+o4GkoRHMaxBRajekEWSL5cKA87AT6D9vUmZwzAG1h0GH8Re
6vrnHmQbNijjIN85PokI0zUmkNLy9WhH6BxXw0LRnZVgCUk1oANaX4fiLrHGs/EbDO1iDskoBVmx
sLH246SLVyioZpgTWbsj5tYvXiwjCcXVozMOXkGSutdglx4mgD6DOrC+g5HHnxPlJy4EekVX/A5Q
yvPd7EmYuAS+Ik3ohNae7A3RTgaxnYHATxgdtfRzQW9Pv4+JA9TrxLxmt6jOt3CuVKQfOiWLoUCv
TU4uJS9oCYMKII3UYR+zmZqmpxL7CNBIre88rFqGo/5zNb8bQrpoMNspEhYLXDTpytAmxyx8Eixx
pGu1X/Jfo1fmYVBPyDmetUl8ig61FYuzQyXCTK4BYxL7jj4+63Z7B+mXrX+iLL/Hser426j6L7ov
/OKFolQC0UPCQn+EEAf3Mg2RJftLe5lH7SOpbxexLt1iTPxa7VwX0AQV7TzOSxjqhfyK/d/Rga4U
E1sqZOCA7ajkYCL4Ef29yXrDZe1wKr/POgWDuBNJtsXTlv/iLn7qxcPi50B1O3ZTP0IcslFFACn7
b/ptYyWK/RJdVqtd0GnW9f4pMHoplN0UWBpphdnwcy0GbFALQb7TpqMSLLvtbmPJVttmuAznPahg
y0LSMV6GrZhE1A4j+Hkg2+8zI6zBd1TD2mX84P1gDByz4M4cCWxuyf8i3fxpWiHnZrawxRr5HGRJ
oqPkkfDKAs4tNnrbVPctRHN2Sj3948en6BaZ5MqrTanxDKNrhyKsV3pY2whLVfTpAzXap//DH3Mo
wuWzfPQ7Rk2paiwvB0ch7PhLI1sDayDlm3jAwRLPDobK6iUxxSF0f1HrVQz7gE0owX8BLe6OwTSh
HnvHxRaLHumgGyXZSUbWaB/Glr8aNIgHjPpZqh4S30Mz03FF93iRD1KyzVflpC1prtTJAFzRfOFJ
EXKDyeta7p54JwAx2gxd0hJYW2RrQc9ZS4pA7tiA1Yq+sE5zE0EdMpD8ytdVCqmbW0jq3YKDiHqp
jsed8bCNI09A4xZJCQNxVwTDvmf7DlKDb2z9NlvsJ54/uEmQI1khf1DIIPu2/FdtK2sbVgaUDD/Z
m0bHvW8ga1sY7BffTBc37p91H0/Ig/AfW8MymWaMN0TzcfPsg40ZrsQ/dRU3GVWvCkb0iWkNqui/
3mEnaKeCtJd0/7hjog+x1ViU3Bs0rjcakLjYdywouBkh6VQTVQqz3sFKA+tEyWDq5GsiI36Kdd/O
9h0fYURp263rpHAEGkce5xrPk3vpbpqBfK+ebZE0wVZP5oW9DBXm0o+13kq5xnjv48vqoSH9YfEj
L1BXC0Uu5X0GogCbuOczTfrAr58+f8IHMQZ4HImmSYaD6LUzApuh3Ngc54YSTvBmAxJMEcUVlfY9
6QSCN3x7pgAat55tro8WisqPwgVtuCSVgLaN8LXfqJHb+8TlzHJMl8BV6boJA74zqWjIkafMdSZx
vK1gM3oe2CxTNKfnhokQFULOMwjxoYNlYdfqWQHI1OeyQbSURGYMnhThUjl6SdHZYVyzp8rvjtpO
avpWDyav+aNhPI/zbUmcGPoc14MGXfbEKthhEkEczBQs8Bq2M6jmrlYWY8zdbFQUTSlFJo3r9YkO
EG+T8y226W5k8Y/xxUzRgpbzEUDZ8l88sviVCSbVxZ4ugygXMCC2Y1VlRUkqmJ2WY8Cw77HahnC2
sZ2HyhcKzoSca48bFr93J1QHCmf6fVgix07Y5cvz/Q/qMFbzFDq6KVx1BbZg0jxOMCfDFrKiDVq2
ngnfPCZSrqJjzKue+yI5iheYekWePV7qTRBDa+NnDOzAcKLME9nvtgG7s6mzz90fHf/U9wb0rHyN
8tXZk5tInLV1xfmreI6Ac8z8WFDi91/OhK0CpMoT2FAG4z5wUU/Z0YBxXZxZjJ6tznvFiSsgi6aB
Rda4t4EYQcyJyu2eVkvKMeITyuQB1jHMkQqmn5x7Y7sCuNrY4QnM1FkHRqQUPYf8EKYOER8wL/Ho
pVehrSqLMtsJ1R+rQk6Gn4qY7q2HAERpmKXfiDiq6XFdB9SDoB+cqBf+u4xY7Z9TXSxWm6GShG1s
XzCPIt13xnaygPT+EzvyH0GNdS3E/FOvl5PmwOpuvghQVwShlfOy/KHmLsqlBsDKqnfpN2E/kv1q
hszmkm6tVR8Q6y40wk144xNEO47utgU8LO0xsA4NAkiKlOvGIZyxc3TrPWcI38mzLNTUuv4pi2kL
QbRwdwetoLHyGbMBRRmAHG1dbvli2kFtT+1bQIczCFrb9wvdmwwacSV8IiRa8B1wTNsT7CPfWVv1
UPdos1JKUp0xh9xvkkmBwaBMEopjLVZZKBDM8LbBHVVy1wxdleOlCRzW62cutEZE7d6NUYWX72cK
umBD0LQrh5yLNdTNXrdGeBh9HvalblXgreZ736JrW0rEKRC2YngfM9NmdZAeNXBMYVILUss+nKrr
fojZAi9gYTv5NN+O1Bq0hgjqK44t/rbNs9BfxNMllKpBPtlBfydEPGFnzNntZ0vvlVnDoWuAYNWr
YB5ee4MAniZH97YrMgDVdvT92Hm2AbD/ujqR8kXwC1kCM2VK2aiX0WHx+mbx27G1+tvjEmms1k5F
NVMwu8VSWxo378P+u5tMfXx8TJZiCRUDumZLn5h8saVInG/ifx6q49pMqb6EN/smCpPirLNAQDVC
pj65gNGd3BdOjLKr/yRDTZIwt6d9wgFawqIFN4a5fCf5KVOlzCpVF72hoKT8h6WuBkRGl7um8mJG
b/9l7QJ8GG6S13ZdSoJOsLUPA0HYODk2HdL7yRNwpAyImFIZ0xsUXt22wa9xWguIDHbGEgTzDuw+
cPWVS6gGbSKmSlk/r/rD0kaihOFWGGRn/d5H4LpyabIiOm/FKgiwwboox4l1BNoaJQQgUfTmOpzW
b3aOcT5SNLlFYbOqgk43vGvDFZk65TKHgAuTYFuvSGZ6mDXpQ/WU/ju7baTzC0KYJWK3KgWbrBFH
s8SLBlDZ8IhTw0bD8tao5Til2DBesykkupN4mpTWIzJnRWY4e9638uU+IJTgi1nVvUoQ89uHGEy6
Ca6NST9hUdnpjr/X9p3GMUt/HgNx5FlOHKulWg7lOFzNBDA88r3dq2CEa9JJpkhEyjNcudM+CLpg
k4xq1zGNzu1PCj+RnR9fuZilaF7shlO0dlpsWmfZZBUgmszhVoGSw4ckzUC5L4Q6sEEmseMkmHop
KNncerEJJyTAGGG8egWrD/lKUqsx7gV7/boUctEqV20/EYVc2W4Aa8kJi7y17BB5u2/woxUj9fr9
GoYvU6cXctJX3aAYhPf0qSup/xwjrT0fFx15A0LM9VV+3sy4vZVSAes6bHhNr1oNMsy4/L7nDwgA
PM0r1unPyaJBHDdapjt7PQMS3gC92am7y+uJGFXl/z7ZQwsEXne2Ij2aSODL/stjDSY+2f94vS/N
/7d9G/V6b87hrJdjFnEBxEeV3aOOUWzfPxN7fWCQTX1YoKlgWsRYWL+4CSHcxe9Bmv+N4Iwu3I26
lkgeVErQehC5TkKRdXCrLjEUAGGh2xaxfb4KfZjLann+T2uy4lW6+971ZSXcRh3XFBo8HlSavA5W
uNVhOI1h6Wa1ZQLsBmVAmkD85RWfYdsePXZ/kBO+gUny3reLaSFCiMjDTop92koCVVQZqDZK0ZcN
ivkyLGuQYPdUDuEMANTnRdcFkWIjREgDwOQ+Mb0BdHyh1yv0LZO4MwFKBEq6zOUPzFMxyuL+zil4
1lo+HjQ/XPaWuACkS0wXVLzakWEHGe9pWoBRgJzA+svxA6CMiST9ZEnA5SgX2T99xXb8NPzoT22A
qT12n/uzxyQwbJmM+Gn88InHm7CDONAOaW2Bjxs0gwC/GYU0QAVzo1AoJS7A7nojPFrqDHFXzTgk
qVjIMeSZ8dx0xKVgA5lLoIOUJxXDlox0K6tbJ3CwejjMtL2k9ICtaisyOEgcu0Xh5pbSqMxoLW7I
/Fi2qCMLeqE0VflI7hQCR9C1AYQZxJRUYvQDuh1CUlzdKbV6m852I1nSALaYbJ3xpS+oPk6AgOXQ
LhjIwaFJsCsjDdl/2MJdatFdC1zOvNeTlBcX2cx9cMXR0vy/VrOWADxMHp7pUA+vjdEaiQZQ47iF
haaONGJCKMzFTTX/NSsfnnfa6/JWlyDYiqPiTfEVvLwPPAW+ueUqlyjtT3f3sfVIQ5HjC6IzokMT
HT/bH3GtJB5KkUd14XR9r7BERr5MvogqD9qyC2TzaXWY2dEW7xTCrprOAEWbyYt1aFM7U46np+cS
frC4iT9xFnENDNk1MD3yPdOgBt3BudqtfwdSP4ndbIV4NXiWT449KllaSyYTeyom2O1dhDW1vqUT
5f9ozRrRPPCbO2W1rRlJ2XeFP+38mtDtwxCQphsX5XiZlcCjdtfxjwVGidQoltg0yOkILmajvQzx
G3bDdN45DWOnWcBLbbUU3Kpd/KGtRLIisPcaJeItJLFESwvLQuxaO+dllV7pDynuGjK4MM382cfX
3kbT6K+9TB3jFuoO55CVPfsYnpe/48gFaMxkNAJs/ucfJPYJ7f2BMHMA6ngFlFDRJnooiH+sbWZe
JJnoiFDEo32ZYGiKzDZeLeyCFfX4FWa8PI3qayYuLA/5eS3HNrLTWkzKgtcEarZsUbIINky2yH/D
wivVxWZTYUD4CmzgARWqkswDo9P5RWJJV2HwqvIajG7BKA96aJPKqxI6zP0Xt1ESGZcjdgGD7mVu
RjNzw5js2ra+0wWXTYdxlHas03sxHTHWy3Rg09HBHqlugE5EaIOGbTSc7VShldQjk1zWqf6jYSIi
6lrt2A8opnNVk8SxRzEqUpF4Nsm5UqLdUg/152Fz0mDOUizG7tiFJ7yIvgeirX1nKR3rOTKdHDwA
dJ1DwVKREvOuI+HbZDFZyABK7u9bujao9FFZKNdPV1cRKK1OAhcePU7w+Te9TnYMHI9mzDpPuDO+
i0jEc7bsYKNX6e8al7UrVS8DH7FDJjX0cfzsgNwA/BtNNYA11Dnzz1ikGvZX+vJIm53jDZFY4hUh
ulLFWHAIVpGBI+BOYSHocMCRVHnOkokSv30bHkOBNcN1WuxcY33mffELIGjusqOE7ZB09ufvj0Zh
P4rlRG/F2e3mhnyIpVmAxQN8u9dCxsoWtKOjCNdoy07YcthAVKyde2T23vnii7iypGgzo5qUGuS3
a5OKEO/CFspyFr7IXRJ5527L8QaITFxajt08+F6iCS7oBQ8z81ick5xmw9/IjWuy2BcSuDjXge4U
VVDNAm8MuRwnv4yIFfLRe4yDBkRPEtsAJJHjLhnKUPQKJmYv47VfnH4rCKaY6aqjnVxbctXJU8ow
65t+HeTwlQvBs/V3BfpN+8n3WPGXKRdbiMyEOoVtYDfDFDErM7eOJhRxkX+aQVB6fuseb2Bv7lVL
6g+jKovivBm4Lsv3sayi/pNsCiBPA2ET/AuakrT78G/DFhyP8UBZM4Vu0fvSrggU4GTq6HLmKSHJ
KMQjTs07gE0ATHiVvPmqvfIvhehu1JTgw/4bfI1m5b8aHOLlGGgo8ogPPXZx2kLnc+D82+pguN+c
//PvD3KM3K+amgtpMpaympKhIcl1qPghDcvaXlvLHSoQ4NUa5c5klkZsWmIVGTOCq6OMGqElB5Of
qIVHsQ3EAkO0yygs3uLWmoSy3uJ88PnbLBN6tIf4Ef/G99EAROLTWp2x1N+3FbKdTssj8QT7VTl5
DTTxGldm0FI6jzhbfBi74DL1Cj2MCMCF2QKZ4evB/+hGrzdghlPqevEEUew1K4umS6dSeXgqzh2w
yPghbW1JKNfUAefKzvMZPgwDZoF/Gg1HjAe5qII7/AGGpbrYVGacBTtRoL/1LJqfrFE56kzpamqp
4MoDNJA/Thf0DDfNgz+V30IOsbJo8LYOa5P4HMWRSK99HX1ReU7/1L8bHZeuOKHi7xYFvrfv75Th
yV+H771ODcEfArb9X7zUj4Ps4D0pWyd8leMh6kVS9XG+VMw8ex33jg4xq7N4+7oa1vEVxVouN765
2tlH2EsZo+rB7PXctF0ELS324s9chnBte88ZtM3ptb3cQTTyDne2mKKJjm5AoAl8O2mEimVtxsQX
H43jW+9PvHicK+nGFQuWu6j6ZqT3HkmaNojxF/wYEbzTMU5FUB/hdBUM92DHrqVAIGG6liVz47A4
f+0wyciFXSLsJF9h2xnuhlWOrln+oJfZppmAPSN1mZYxdGH2ZDYLqYplAK+RP7nmsBZAGDumhYj3
vAPP0VEIcu4zdCJdmJ9DZdAYzR/sQ+Ibi/XKM0CzuasRGCOVhUiGS3v7E6Q1KmJrAV6zYWg1Tf1v
204vzgP96KUtD1ki7ctSeSkN3j+nVj6UqPvITLhP7BxH4CE5GR5vKZN1YXuE1IisCszAoVR/PFwS
aU9NwtTKbD13UFa6M7oDwErqTGd1YRWOwUUqME9wsx+316ytPol9b3dDYyemiHbnPID0i8EjhOGb
da+P2vrK1YlJthIryruAPzZokYOXSpiyR2dhkeGp+Kr2JaE8IVv7dtxhqX/7w0KZ4jBnclh0P5mY
ga8pjMhwP569ZK6A6ITnR09czfZ91zBnb1g+VRMJPEmu9JW8MuvN4ALkunkoBP3ot7Vnb4fi7ImZ
k5sFBYbLLKWAMCmx8TPZ5SW0+4LzAgR82Fr8Ncn1LSt8CWQ8f3qfFA7uMQQ3S1Dd7WItuoi9GaRW
QGtoYom4bf17uARIhDpCSOsc6i0AsvUKGVq88tK7YGkTuNFLMaobj7agOWo6NtcbIfEI5x73SwEa
k+5yyZuJA+qMq1+FsCB1JvaWST72sqEcJEdg/SwruA0nNefvQ7yxviIfc3oImY3FM6Mboq8oyqkk
q71FBAQhd2rIbfXHG8DnlitxQbCtulhP24AFsRQALDd814VZqUM90pUX5dh7fY7f7fnvGM0S83lq
TJFNAQ1xjgodAAxOsHB8NUgLK1emL0X90hgpZ2OVDXFm2EPQDQTs0dLh5bhkaTVKBQBfRC7PR/tV
Bak1PSKgQELZfceod/v9F0wVdqhpq86W6DhP3SFEvRc=
`protect end_protected
