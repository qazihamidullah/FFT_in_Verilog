-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ElBUH76XXt/hEROT3ioxr8P+31isFCdYmWAhl+Flhr1HdmAhjXIxJ5xfvwVVpTWFIMZytbM9OXoB
kXJ56cSc/0YTz0mCiPqCjF7RFjpjqIAmZf/r6sAnFrHJU6mtu8gAFRijFDc6uv+TqOOAxNzoLNzK
8c3kmUVGrulWCO8g+Yskfr4Y0hQYeV2H/uy3jC3pqliL8kvC9IqzESt1V67WT08gD4+yqQuPUr5L
yl41xSkITjrWeg2FDodf9pRXvDsZvW168QovUK7G0+CVNL9NPofNym7hNg31m5pwTDK/kTh7oDO6
k4GouguIdos7kx0rVd+PFvC8IK7bLaK77ZMu4A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12384)
`protect data_block
ImymGZD1BpV0A+45Kc2axwIuxef8qldFQGnp2IGEOo+zYkAIegYV20h/+KDjKOdKkk78J297ZgyP
O/ib0jVqYQdHtnfNNiG/MF33mtBeHbZKMPN53GorxWKaRO4HwMQDTG+JwRJ2ASo6P8Ip1TM5qyhf
Y2KNtATN1XNoRgC9OsKs/OgUJ5Q4vNICqEU6ltTfR3TDcbIp21ThkotuanVFN63tt7KFEeDHXxRb
Z5byi7ZcKfKZrU52n/4DToITrpbhlDkOVk+1bVWYcqKcwvGpGXKcThDeeqJuvZb6Vi1df4v3R+w8
vwrGl8KllZwLHBAoCQzZBDNvANHiHZ6UU/PchjY3PPh/+P8YokWZcYS83VN7fStlnvXxG4X7YTGF
2SjBcFLMeLD+dwU7zUcD9Ir1dCEJOD+iiO/fJjxHfw3xX7Dy2dVv1dbHaanGmoo2/lV0pHMLpRH/
Nnclsvh9WiEvowtIjows7FQJkY3+wJhqR/j5aK+elwIbX632GI6sv1Bt3+bSbfKaPoUebB+bbW1S
L830GeOiQCgHENTC8IU0KdeLFG7T9erriEdhNvEpJ7+kslz3lqtgYoVdW9og7imTSDbbpxMxXZIH
ww6MQPTeTLv9GG2En/h+9dAR10H+ZmAJhwafEs6Ii+1nx4Yy4TL0RtXZAMJCmp2d2nX8ryr2D5LN
GbohJ8n1NAC/bN3X7QX89GGNwG4pGnfzx3fFaO6z1IuzI+sKPW7hEAtlfJ1d8X9PKwRjGLfSwjE3
BTkZt9oe5EWEyAa13Z9Jh2pML50LCMJCaLaYqQ5ugDPDEOH4NJ4t3GikIhHxlSBtR/FdRzftDw2g
teBz9rA83Ca47I6PNz9mQMFjnof4Gy0J8XegSz9r59N+xU2iBRKlQWN//1zi9Pk6IdogfiPuJ1CR
loMSJ6IhcsJfpNzSbqXEqHk0WcFW3zOL+BDFi2Mjs6Du1T6+MyNb2O8wSbcwkFQU3FeOeGJ9h939
oOkUAKsX3HXtPH9Qd8byrjn1fJsbVCIfxs+YXkOVbHTC9k/Xj/nTaJh18VZbHf2TSZBRnoqFbuKh
d4YKpTYVv7hLo8Uth70yWsv7iyC6jvBlVL5oR6nwHuuS+kuzr4yY7JP+knMqLBBVdXhFWtG0xagC
rsFEQnvhkLWlwBoaRkEoKQErITRELjKmQYlnVK7mF9lU8lb4u1OnYQD/4bM2DmdNUm54L3oBMqRL
aFsSXFHYlKbVHNs0lTHcCFV0t9zFjtFbDIUAWcMdlpxZq/GoYCchjtUL5eTcxCD6UunVSHz/zc9E
caFQX6T4b3/g8btmqEvU4CLxTjVnYr0BdMxtZiZT/YVZcLDqNBDA7ouP65k50TfIN1pdR0xCl+T2
L1CKFwgeLquDZgRK/tsZcpi73f79SIShWZ9zAM/o0Hl+m1u7E039KELP6gj8rFamJS2b24Q+EJNI
nZR/Pwun2P2JfY8i/iJMKcF5JDwFcHHZyT/1/ySOlDGil/QokeOK6cvNyoG+5RsgUgTKkl1VfFkm
r6XVU1zsWKSxQ5zNiNzZMyhsSAVY/Mc+bOmcwLrEZESeeog10mIRcTvV9tPsf56BJ6fDl8fMHJC7
p8pXu1uOJW3kaQC2iOruWXrneurgrR9gwJSzkStPUd4FU/92NqI1JVPxy01gPw7BhiexK4qNwzEA
qjp4DAXmWZiV4ieKBc95EhwBch2cNLpYwch56gYabbJlRROMLAkOyiV5d8yAJex5ZBNRwGW5AThY
QazEQQzxF+H4qIgN85/O20qipcbfQuiIBvJxhKyCd0qByUeQRSP+WsYTsJ17/6m/Zq7/FeV8kGwq
mOoe1t+Zs8W0+QFhrvEiS+URyi5AEFrPDkXMII+Wgv9qliiBdjjRgFIflNfQObAyhQl9lFYdiT8r
3BqTsm6OBXVZyg3blF7Hlzbk0Cv2rGEMZlwOcqeY+YqlMHkzFZB3RZZQ2ZR7zrgDFf3L2El5F9pK
S+IhjibiQhPdvktD5yDAs5uq3tA2bgY/4GIJj0vdkXygRlt4XyD4GasF8IGDj/ArDqbW5fliIDHR
PzYEnvyMGeEP3PLeViy0pHgnVcYB1xWC+yhE/vOBgYM1LLU2ratXxJYfhbibLlVmaYAczl5VIaIQ
a6ywO+H1lZPkR38lNQYM9nUBasABWCjjDmJduIQv7b3FkEvat9ijfCXQLDM2DyKuri+tfzqwB8CW
QRx0wgYoATW6sX3k/0vcJeYuvshUeY29AS3AqusDSo287YF+IZ8HJ8mQxAw5E+YDNbnla0f4Rc0F
rxqixFV+emJlb5EcyERr/OsSPeGkAphChuTxOX1xPmpD3Ry+/O384Gvcvut/USVVvr169max9noB
tsolnLl9Uo1txPhh2gXwCDELsob58Em+buAA7sKa6KTJNTylbE+D0R796lkZzJlLOv843t9F4ae8
biGe4KQ0zRd03gRSn/sDMrdspChLmdIhlLY3M4xgsajyLHgSBUcz+u+ovSR22jcKoh+5aHUq8Nc/
Ac20viha5O1VIotctvCJNloNa7dytAWUOY3KSNt2maUfVqCP11WtHNnbFikY3uKHLz7e0Et1EXeU
a6tV1vYlRvChiUUPgG1fpjAZwqibjdIPXuEStkYhxtz22eTkmeReWGhWuILjnlNRhQcmuszVmTyM
4Ew3w/OVPbWHCLunWs4kDJn/ggoJ35AqaWDP3kDvIcaxf+OndqzPbcOdojPZxnM7U5J1924kP20d
Bw3+XyNXICkQSLsuqZMjzhAR5btFFetYJQgDnN64Yoqzbo6r1j69rOefoYq6p09B+xH7ZG80eOwa
bYeLczu0FSXa7kaghYFOFV1x6kMasuiYV6I+PRNpgEGkDX8ZMM1TSa9KcMeuPUNLiFgdXjRcx6Gh
SwEx5ENS1NRo/dDPLtS1/lpAP7sneyhVH/e+dFUNKHY1jb9JENTyvZLYzl4Oc3wCcQwVGPmmXP/G
hiQP5aAsOAEQBJNA5GEGIeWTU6mcw9OUFuh1xWTBUoIhIU0tgA8p+H519Npfrt13D5krtzeaDxWj
Nt5AMfnE+EtvWz07irwkqb687xh+mYKHzqdl4A24j+WkLSu88weoNi8+utHJGO5ilg4PtNWiWeu3
ZKuG/ofoQpW0k2bbuJO39zY76A6Ym5J4zLIkR/aX5uu9NiEekaajBVisWSQjwZgnDr2QCmuhMshT
IzFSmiqhMOVLn4gqY5WPfsI5HlXfi/g/He3XuChCaa6zrgnSIllpdW8URhvfiUnIBeBo0JOAU+v7
usm1EO72ZFOJcWwcsx///Do7D3zDtEPTD6IiLXCd8737YGafLFw33YGGm6kLqUSEsOBTKLVWUSs1
gXviNga8dgm3uAnO2ewLcxiotQyVNKFI6KeAj2HA6aracGekIeC8VFv1wkkF83nCmMz0aRtdyHEF
HPnbVX9PmTsi6QfY0+zfOUFZncpt2tS0P8wjdCm3o3X2dz+a5bOkl1l03iR2qpGh0BbhbAEkNdvl
mNEW0vyAktHFPE3yBe1ruwY/vlLudfU1tBWpyN6Y69+WAl24gFkh4gQeESZs7iv9wbIFskwjZtnu
P+eOijcPxKNhfPYW7hq5/7D3k3fa0sydC+0bXZ6FWD5wUrkAtrbyvLs8L0qfiHQaZ06sETuI0nWA
OFiTG4JZFhi8miqMl6RQvu/gv97Zvt0yWaGeruagzCRdQ8ukYj1KMpgnsEn5rvKbiAKQ73VHm5Iz
rdl7uJrKu+NsfJ8vlJv/QIHSnZBQSO8DpJ/TWDW/XApjvkzFzhYoOp8YG0nIIk+GWd3shxguzh8f
wCoIOZ7KVTTfP+Wp+IbMhQnBK4mNDoHTNXTtZIUrKhReluXNq5J+3mUQdJQRTv8XYN3quri6BDnZ
OeDg1YiElpVAogzsYnuw6bfr936ULdCFaFmSuuOjr24R0vZbMVFtLXXcEo/l8y7BkSy9f4eG7Qmr
j581jVp5eyGs7vyMiUP31OtMDsoJtYImwnRZLow1+3zw5xnn13qI8fNGGTXkBq9+lyd2ne0eVMzG
d0z0zY/fiz8xgHQW/5ckAu0EEPmfgiER6wr/0Mv6FjlVMu1Vsjl6bGLS+jHPVYtwVx2KlpPJUAwV
XEez3qjF+rVnwGruoulnGxCuEMJ5aMG/OT84dybkPszr3/IFTS5TQv5w/xEwvTA0x4OTP1CuePmy
+0mLAM26mBoU5UdD68IefgZ6h/HJHGS8jiaPDSraa1xB/urVAUcfi6ZeuwrG3mFqIoUWocOm+t+u
S5T9VEqZTrFxUfAxG7Z2SWyxtIgKA5zHyua8oOPIIgMoagJ4oMHQDqJvEj96J9cTBtrdFYeIskGZ
whokmUIMfcmXHi8SEwirSpZa5qsshf5/zu+nGKdTrfLDL1Ce4V9xmnnfYc8ZVZdVRa0+P79MT+Ip
BKQG5z2cTz5KO3hiSjocEIb0iWi0q736vC9Gt5jgLj/gEELL+PY9XlS5qUbqLNXQxIrBA54WjQXX
OTcgQkbtliZcgQwgMNvlQiJaUQ1cokdIW0xHARox+dHV+t6LHWDEWny50u6PBQxXPE09aqXs/wze
c9GbsMVkH/tPCW0c1cXQYQ9yyWmSF99atAx2a4DtOe7Aaz+eFArLsPLtchhAjzJlqbT1O/KrJPd/
D4AZfu4uI8l4W8C+H/OSO7hu33yJkbfD2XSW6EDzkxjnHAhMsUDQ3jZZiRyO4OhVPC/fAA6J505v
uN5cr+VvpW2MP/o5cRnB6VdfMmtKLe+f07ew5z7I24p8flHjOh1nLRcWEPzUTTJAalwxb3sAPp/s
E8+9wTvMiqUhqkgN/Aj40scQFxre59kPP+W16zpExRhrlCdNvx7jszWlNHIMWDGUSrR/yUeCpVGM
BHt/h4BNGbB/VqJpE5TFHQH4dgQ3sNhpukxm8YcQJhRTb4GKeeiLgK4TrFrY8aqC25S36/7CZ9RZ
gFydkevSQE4vhvsY7kaRM1d8GD2D9EZxpp5yLZPacxrcLqqcCXrDZUeOQ5/XUuAFjsZ+iFdNH/4G
6hECXE/R0yhtfUU5FM3vKilU+bYVgAcLPLnbQDSFRsNJJvvCzuJBRsflhqURE860h+tRAorF+cQv
l2UnswxUMkxI3f3hdzoAxdz2CoNkLuAldKHj/TYChgotsap0gdsc+vdtIbEl8PpjpzFzW2OW7TSI
6S7LSzOHicTQ77dd1/dNgYDToVJCs3KqqxNtEgDFwtO4WATX1Nuh5IbNCDPdlAcdHvyP0f2pPjlt
4WzO+QJNBLquHpxXquaizQ4YotDwOBcGTwZkJ5KsdU8x3jQGvhEp1rEZy01X+j0gp7C5MEKV3Pvn
J/gwHSuY9uCLqLcCQrC3AwmOmVYjeweVMEm9KxDChZmc8GCtliasilCHjyk8zEawtdFN0Ag+E1wU
NUy87zyWn+pUKG4sAkoXs35J9Qp/h7AmtpGHufZR2vGN9zMRHLgz+7zAt7boHTjM7zYuwWYurMjo
RO9h6mz6kcZg83A/e3hLpv7jxyQNYNQW9G+cMSr4M0Rsd+lf6pHl91SFi/GvYDHYvyXd74+2n8us
BleR8/M1hkI78U61OcHu5WdWiqEUoXRvUuQc0YRT+oaGAdKp2EKucmGHfqt2n+67xfrVqcoaeCg6
uy+OeoV3gmlHV9LFwdbHDtGpw7X1k1Rws3CVyDT3dGNwo7rzLTGgTODXTJKMphaDIsdhzOFQz8C0
aryeDlU7868ASH6qZjBfG4GddBi2Q6MIsPdLwIhlJqDSlbhniuq89YEYTcrRqLKCIJEyf0qOadFe
0D4Y+AwnD2I4J8GJ9gcE8G+/AsEVJ3AZiz1wOryhUDdZcPHWCVZnq1HCBXnmoUoG9YebrjErda36
AZy790FKTJ5CXb6a+VMWTWYFfBH/ylRg8aApw+M7R3y74zZMZh9FFXwYO/zrL8A4VWC3NpBkc8JT
NU8iT7OHL++nBUGacnWjyM2vvLSTNQMBQ7a2fHhk2B+V9yK+oe59i3IpkWTm6xNRQgjAFZ7JNyxx
7n3hEeJ85Ji4Bw92LnMKMAoFS//lh2KbZGR7cuvyj63Y985w5pbr159v6Y250ETrnEvEcA0WiJTL
BMVUnyN/o0XG9tzfltaCeEoIgFH9WFBKJatGDVkaYrq8NvRdMPFg/2lQnIM4hXxTHyHyHc7tKyeq
T9W85lbqSNgbtmOY0wDDhKfjonEoGWpekPicBlDzhRzPISOoftX5zw+ZlSvwoqP68mfQ+zX8sg+F
3LnCTajqgXiG2NY9ZHjLM0SS/cFpyPvhvAR2HZ/YdaUwRnEG/YRVkHr1+Y1IBML4cHCNxsP3DYp0
XFJHTA2mIysmPdH0jS/LCqUtdUqOC+cfE6GbIOXhqH6jVMcbQP/rPP11sEKFt4wRFnYnGbkoCqgK
3cPhXmPyr1yJuGLqH1MmT/jmcXgy0fGQYzrwaGai5ExAMMjgXd+Ok7OYFwRSyYG36ygtmSYV99FP
NkIJrkSlQpiUtkFxkwBCqcqZ+2FztR1qEC81BPaTKCvk5WBaO5kMgYqi/uHfA61g2dUWFrYnx8RD
4JXUaS3gvO3UYRB/8mYjA8bUqrr6oy0Ns3KnHngz8jDDLEHQ1e5ON0bZvthQGBvVs2D6cZGvkPbf
JeZ+1aaJ+PujfPZoJM8hMuHW9fITPvKPRweNpz7Sg9CGTf9NeLMOP5ujkHW08q1b+1cpHI0K23nD
Qa9xQG8PnsedjrGzAYHov8th8jAVa2KXubvZB4d9YwP1h1v4x6NdZq81ROChgyfmNrNjWfyrQNOj
wFfRYgPQgVXS0K04roTPuJFBItd5AIYVTHC7rFthCYWi7K/P+9eeAnfW1Hn0RcpHLv8jQ9HRwIRe
iT3wJwpZc22vYZI3/kwhXulf0KySeXi6nQm/H50iGsO1WpIe+cD9uBoG6HYgpSq9dR0YlLt8fV0R
3oB4jHsYBoKBaVyPaLoMUxSDnQAVqeml20Z9ymrxHfYMgb1fv0yrF/17PHZtSM+DSZEVsygGbJML
G3XYg5tLTa5EY0jVjmFWieRW0sIclRTjntxhHJFSikyp1+3QW2S6oKDGfVxFv8Rk2qIvoOI78svO
Zl9ZDiBAubQH19wbGW6K8zlwoEBlm1A2ZtpH1odbCVBFX0XpblZ90RgQFLZd5MY8xNDH7Hy9iK/j
9dEu3LXEgtKdYQKLHsi07ALFCIel3l1NWS8uqvxo1mJcmz+5BtLNTa0GRwbkncDJ6PF77gFK9ruu
gTSnU+j/YTqDrHHKhE/kHX/qCwfOQTmNaxqXC1t/MLXWuR1oJ//Pd7qkacNgx4kjoQPGotPx4KhW
K9zaIh/gsRDYefYnZDIySg0TLiLbk4/g94r+SiyS2jnWvsmFH4lZ62DCpUx1l/GRtbySMZrPmPRU
9V6IohCwMQYKZjWIQKANlSql2t8wwKOvWo0mNI5CjwP+KB0WAIc4/Wu2RCGeTgutNgY1hfk08mHp
0qmaKfX3nZbln89G8uAC0oC5VqbqhwBU2N8rS8CRWnxcNzdONETJB/uYWIOuItKLaU6AgF72YqIb
pDScF35ZaOjZFoa8HkzTU361Rtb5FeAeKM2WP2yL33W9RGo/+Mrn4zJSGhj1R4lpbtOar2DlIVJf
omfSgBVvRx8DpsTtJTJ+ttVKWzbUB3W8kWM9sGz3t9pjTSQ3Tw3tF7md+pjc1XdC2i+iJKqQCee5
YZ65YgEUBQlwF1usRTsyrdpYsDVT3a2WP9b8hplV/TYMfSvOtax+WUV9S7aDF3SL99dYzpHQvGJA
rV1U3nIL0LjYFRwyzWxP7I1MiFW+vcdpLDVQFaR5P2VglLrmAcI68JtV/LX1gjKv7ADEkzLngUiq
vZzYDmlbLWHDlXyTi7jiA9RVjyn3DB2O6M4KhBCeUerJg8yloI5L/xY1fA/2rI9zcKK2D2x5EMAT
Om54V4XAI5Xhpj6B/ZHXlJt+M4Lrsc2sVIOlAIKQbV7XhK/rWwxX1+dQIbwOuV/L2fFJ4ZJUxtxZ
OMmCePqZ7SnXPIr3HhQauLb65qv7BA0zhFW3i9iSOmVr2QrshgKLM8B78ct/Tm6iRjCiKwzG7tcx
LcbqO77DmUUYG0PWCT/ODo94WqKfgUDxHreojtOEXwC3YuXMEsWsBgmWzo+FzLvi6gdJJiZ8HQr2
/aIJ/fxQXg2LIvVC5iiHuZjUFPAiLPFCH7qc78ueZIw/4e0zP8+3iDxTMv/s4iShWuTkzI77GOm/
p8jiUuz5iZSgOoxU+5mhh/xUFSWo6h8pcQDVnDaFmnwmMm8SNtG9MYc6sNPaeUDM+z3tDgST24ry
c13bQOPNdW1NW2OtUmUC00C50pqEkUTqAL7MHxa3j5I3FpNIKiAkZSJAqA0d/7CLHaQZbz1PzQz2
fyogthDHGux+EE3xgqYHp/JFW1aa19uBNEoMiAn3dRgrO6bMV67NvKAR1HWn9GzJQ3B4u2kRM/qj
AUyIStodqRkF4a6NCXVdwjGdatTu8NvSL1uTkDrcKkpZXEdzSTv4mz/Jy1HOS6GqD+A6Z7av+wJL
602z/O0hpzxIwcrt7A5rNuHh7q43vFREK2iei5TOHvxkBleh3b6wQbxOyJc1y2vpQRnwy06Zcder
5oX3WBIcWQiStsz5lg80BshUZ3HT8MDcxizM8we9uNYBNmfrINjmT1NHFzf/Pbm1tqcXTd0mS/u5
nI/Ov3cwwIUt9NiwOWJmiWzCplfksp265bJcl8Vr6UT/IqQQS8M/Meh4x2RwSbr0oHy6iCCyJh0p
aytca8MK7L1VKRdR0hPNkMwFE7cqs7Aez8459sy2t/sHrOH0IzyJ3ktvbJoq0UcrxIuEZptaVWH2
zDcGS0Uws4MNh3Bj1PdFWxtSqQiukURpwoeelQRTQ67U40SaD/m9nPxR5hrovTcop9Gkr+SbsRgg
Fx9hqQ++HD7WM8mmMPDY9w77XvoD28e7xwIX/0yC0ZeuDk8se5Ow1YsK/SxNIW6u6srBg+etlqKp
581r5gbCbjAmAUj75iuqzgL8Bi31YV1aSecZdw40zqQotk8Ao9UebubgOybI3ErG769wzyxLPYFg
AnfuDxYaZFPVCRYW4/4YPXHZB6EQIzA9RiMWywCf7B4Q38Cpnj2RynLZ4k67d2gObhD4eOn6XRHJ
HnlUDi9vJXCv5jQIROtCrtOEJrBEFHFNOBgc7wMD/xXhrq68Z/1G/D1OKrih6Qe0e0N46O9DLDD/
4X2wzzS4CcxYk0yIvgw5MVfoyk0ZbJU9qFhAyCvgSCLvlpRNNKtKo1+PJg56w+iehhWVfkOmKlos
DYreeFen3JYTL1UrIkKQbQ724EP7BGcABZEMj8MowkGe0OHkFtUzzfYOVUPY+xxXVKgLjTD7cLW1
NqnBGZ3uDsCa4bynLDnMCkJk/spDyetRja6RNZ6rKLVwveFvNpdzoL96WSfIDFZtWWFzSrQsMII4
rPihBD6Q5rm8c3+bxxa37byS/yj4OiM+swu4T+DyJlN3jIqcUeroP/a+43MnZaBLLlPpWCDiYu/M
tmd9+86sddm4vbUiC7sLTNbSqih4q7wsT6m3UnXoGHUxoOby50Rh+l+Act2h/hJTpsVojuA/cm9T
Ug1yPtME2IQ4EIjfSvE5SOBDcWi0eDhzh6gD1TSYjin6Aft1lNsSCgX7D94U2hLvQPAQ1LrSi0+J
Y9eSKHBH/9qwMwTqaznaI2v/p7AyvQvPUemkroNEwiTptlQSB4ffVm2P/Nsk7vN1GqoA4TcJPFJX
9UqPlJKr/fRVu5qGeoWdGcEK8rhQU7gIpvbeGcEDKcIBGQ86iT/4GDGo8r24F0BftTT4m1diVLFD
M+6kb1739NyTZQgw2JxWhWEcTnKn9ki17roxt9ME/6xwBXcPNX1fbH6rc+NkBGR34qUoZzHnp6fS
qGMnOZEn8qNV6Di9Dakt4QCfcKA86OgbQ49zww+/ZTTqLZdgTOSz5BcIHsgWp9kuxd9ul9gvaLRu
itogT3KPgTRAYEJC8H+RSVUdIf6ZU8ssLjx7m5AG7WB+zw4ykH5nJPus5/zv6nBgKWatiWXRARjE
6q76kYPBgcLtMTFp1nRI8zpjFboewQHvJPITaGDDLjHBwbaS77PToh5uUDC5pKzBp1nHDo+iXxPC
awj04Kh6w1KbY+rF618VPdw9WpoKQShtfC5IbrKD485Ln+7bcaXyCn7GFeJ4UpLtj5KVpyl0fMMp
Tm6NQfg1h4l6IAIlLqPmUSAPw9SDxxomjn3Yp0hLv1cGv5FdBzwGK6HHRZD0hZoxw4iiXUpc//yj
8MNYTLa8iIZD9igGN9ZlMk3PFwwrBZE9HiM96DbFnh32ycHhACDJ7Atwn5af386RwbdDj7GhGi7d
dCj539ChDmxdBoP1kaiMG7qORgJCPpKVNKEm6Dd6WTsgp99EP27AWKhviQIS1EmrBIfHUO6ZJUF0
b4P2Lye/f3Yx/tX6RCWI+JU/zcA2zB3p0eVSL1BKE4tDoMiSp4HM2cDXjZveyAaWe9MOFpjOUQlp
8a93SdL7DM3X+8U5JixjWNKAhjo2J3pPkk4sdKXhUbzlC6Sg6d4eUeZ8cyIrZahJChSKa/04UJG4
wkujbsaOf7zZ7k237BKpjtrE4Rg3p5yEvGJLJbnA6pJqYAvn3jErid0ZH/gVElY2iV7YUIFhtaw/
9Zd0fnFAmyXP+xt2tb63omB0Awbbl4iHbLOGdsIRBXwRX97QyBIMOEeQSMRv0jCVjmzTmMcNbRHD
JB+e6HkJ+DNLpJITNrVpzOziWtR6a98z3Eg83tOhtuPJLq+i+cTmiCy/YJKFQwjK3Tzy6gGcxTWg
gjUrnWzLxF0DBWIooq8H/Y9KntdA1VzJNnOX9f3rDFXk3QKdVTJgnBo6mYUp19+KsU8o0z8A7Fr+
yypy+O1dPpqmcCADvL48VoJYSJeZe5MHuU6R9oJfDiV8bIUSZ+9erB5Pw2m3v6wLVnIdoEa/Qzye
LDujAlpKgUuuvDXvsd06umfbx8kjeeP3S5+alIjFmczMFQQE18w8trZcKavgetzINM+MjnCtyAr2
3jCzs1Av6ADDXzLJvtSfEJIzT5uuw2Ac21N852Htrv0oujRAdd9b3CzPF/knspYvRsmM4WUYhrK9
55uVwiBL3rrzyX11kfNTUN4o9IEacxOmHS5j0TFp15vENa3PZwcqyi+f4pf3EAIkX32Lh75wdQHF
2qXEptL29dw0GVoMsZqbrv615ByqRyYxpXhhNQS3zUAVgH3e1WNNAN5/27KiOrMZmc9U9KFn8ZLz
qffbs/giIgm3yI5R6wvrFC9TE131VOeqV+7jKCr0lHNzy3Q3nmOSV4ZjJyIxc5HykY/NBlKj4K1s
+9ySJQu3ew1fLcSAZF0iPvg8MQOSTLdHq+b+3EfQFq+NdbLAOEvD0lWOkt2tJVLy9S6gD6b5TdAF
LhSYVOdvxo61uwS9LMJfJXYTESEaGav80MJ74EfKqZgl7VxKLveShKVcSzgNjPSZCbs/yP2+BaoV
b46Jigypnue3uJw/YNjw3yZPysdz4HV8NGramTi0y/js7q6a+WDh8p7ZRfmS1h3N2w7ET2FBXs/X
Bb0XVY3fthBVfzpbmcaDqXTLMX70W8Fa6GvmlAMGRpMGcRvGB5hiEwTShw995H7NUqZfwCV8ZxAs
iFl7x/1pM6HaT7jxi6hRYL6y6nfLNQfmLxhjzeubIroZ1sJKmqz+d5c/MlLgXIqTJ71pCS7+X2dl
zBcVywMYjxwxYYMGgXLtwn1i4d/OYVj8uW5ZPIVu8EzSpLEHsHQELG91P4gKsXFnrLiPWo9bOmC8
kCJ6wBxl/5zZ0GYMHHY1RZnbCPrxeNX7SDnjCrPunSaeB9l+NCfqMc1QY/fsrqMxxmvUxaqTwZlN
x5GC6+8emUz2wxnq0XcktzyLDlkupJXb6CvbonZQuzumSyBs+mIez7epTss9QS+ljuljIf9hgcj5
xxfJbZJXjFmhn+Vn4GTvFjHe1trdN5N6kyIOU/swIcaEquIax3bdO7pwctcJrKhpS/O9mzC463ha
oCWHKRdGSBLaRMbG9hQNtMEQEpaMMqoykSylcrrZh1uthU6lzxekk/0IF15p2i7mdk9GMFN2LFKS
6Df7DJ/Fdwarh2US3Sgk6fEkFSuNU2DzcEnQcZyAeIc3v1A8zgKTDLwjfWvKCY88caODaY0Mc1T/
jVaE5Mq+AM4wwtLOZt3h2QpK0Da/mu+kiBuJ4+YgoggIDTvGt068noOP7i70xjoScPGMRfmA/g19
X2DIZ/fKAYxGhOwtCPCY0O1Uvm0Q3pnWNp39P7hMGSOY2Uk9TYwitPd+DrZ/tantuRoSzhc5tUcp
K9+WSengS3bRWkYBc1wV88aL3MvEPXyB6xFkVOkLh1SKyr3lLdNk7voTOAIKAQP6lKnJcGt+V/J1
2YGyTrI8YsngsSUgRB7yKLG7cG9MZ2o6SFfWpTKXENNhVZthCHHnp7a6tvGX3sVaYEAS6Pr0wFaG
9KkcZoGkGY1U1dOTrWTw7LQ2V2NJNWL/JrKvI/Ur0bq6GGl3RIlwKgrY2oRzoLyBlSmojY19nqgo
qRxQuS7pj2bWyAQD1ydQQU4Ay7HQvoISkeVAZpsln860tqmq1q6A0gjjLeo+Lpln0bOgH0qnQsHE
WPoia7jEmIP776Cd/BzOPpa71cjdNXG9eIZQnct/vBzyokOek8viX9j9/00QDBVZ/6DSQiUHpSOT
Y/B5J96qZX0fRgaOPN5pra37wVYUjjKCEQFr6PmSMo47YZLTrDh8j2iNm0i6ikK/j6QYXYlRddPL
EgSbHEe0gz/ZXDq2W83Tdwuvzum+p3IddYZZvilbJOe/J1pNJzJyOw0nq/H2yQtiMpeCp5ehIuRf
ipVC8GdG9RY1em2vwRtEqpf3JnyGEehlxZqudfToOrREAvqPVSQMqMZFeBhYteo1qcTnteC9CxKj
4ipfgJtHo0bPvvk2CA/DuUhziuXzoNqBuZpOxIlCY9RRfqUjAuC7OevH3E9t6s3Cjs+/CCUb0Wh8
fIZCbv7yP331GboAooD9BKzRgvxfRpzrpmasSqf+33qWS05VhZrzKZJ/qOeKoJT1TO2LIRkSAYN8
D8kCkuOn9wEZ7YhXpOvwl1jNwj0hC+rN9YjIwc3hKZwN+oCiap1LSWeWx3wwvndyVEhL8JnAuKQE
tHl3ThIyvRatr5rxRkiSccbTDNGORUJ4HjljOu/mGEP94hXazEvIpRBNDC8kjSyal86gs2G1Tny3
DR3bzOY5H1H8iOKHPtT4QVGUDwiN1aCzkE5Qbo2X6xtJmSojw8LRVO07FX120bu4HcVxTN9EZYr5
eIrNTZ73AL7mtiQFBlbIIyvRkWNgRPnHPEETIOg0Caqw0mlqmny5RuGgCiJovg/B9EibJ7p6YPbD
TWvADs/k15PV+RL6gOGq+eZnhAslvSHPDqJ4Sc2FfcbMG+WBBh81dvCInVcYCGiUNLjeoffoQlfG
edyOQCIEUU/bOi9yQgkfgOmPALPIQsYMJx8OwYeJvArRAVUXrhqkMLCtYVtILO631WlXuoyDU6HT
3TdtpOT6zG0KubSIdeur0jSSqTSbCUyFioSwZiRbL5WkpbXig9fparNUhEqM0zMuVNSS/ptJyi2G
ibdzwfJdEiv/ZB2FUnYRWgqkse1Ml6X2Byfd3s3pQ8bk5jrWbQ57PPZIh5x5XZ2lo1EgkHtqvNR3
wHG+IBm23ZaoEL9uIXd//CqjA9oTaKHObI1acHhMzF2RYLEKLTflXjUtRowTI2CRon3D/VtVBHtA
nOAz6YVY+iPD4PMADd52pPf/8oab3YVzeKclbykOsLvfvzQyW6d+quMPEo6rxiugI3k+v/0RPv2J
1KeEAZaH3Xlr8D8y0WAy7SNa40GYE8p40zD6IW+jfhRuglKo8jcvci395d47gKxiFrl3BO4S+ZHm
eclCwoKCUQhxaylnZZw8u4bXwdyuH8y2g/ikt99x4WkmYj2953RvwStaHlWIewPGVk9j4NLsPbl+
Anjbx5Q3UzrVkHGQT1hfSOVvz7Dh3ClyeSEWvHRbodQH1kDjNvPeZeqzSC6kqlBoxC3uhl00AM4Q
wIzst/9hUk+4RwanY3RbrraPaQgcTR6jvCMtg50ySXHbwOXRZQWSrdTC84Pqu0WNfyPtINfbkbgW
i5jdjL61OKGMBufd4VaOB/+z9Iv0YEu5dPDd3aR2wkpn6fFdefgTxPzB8qZRtfsrmnqeulFxx3IM
lkQujH1oa0d6ihr2gBg60XIjtJDu+x4fVMg/FhP6IHwPg5+IVp+xpblMgTumHfXi53ncPSZRmUJu
Wj4Dphf3HxD3NekLYNcHTNBNHY3i5RJAJQNyDeLBE/i9LCFti+ri4KwwXrCDVBLrFCK6btCrGlIY
nKs0F6dYYHc17GH3jtbcaA1lu7wTerNQlq5omAOpo/gv3x7akBcp4Rp1d0vejE4cQtqSynrHGp00
44FmvNeIMxvDRqv08TdbGJk9c8U/DbMeXQpGiWbCI3yWAmZY6M212aBS6i1kt0SbFelQrjMKoKOS
WLhvPo6TkghfipHZNWUSqNfISXxU3gLJL72G7yE3azt/7T8K29aLmCgNa7Ks1Rt3mglpvStEOw2H
GYThdFSIh2YVCvX/Uy414xxWR/atgKKWon1DADMqkvr2M/CMDQGLJ81MPULdEt67KxUA4kMfqP/u
gd9U/SYzhiLQelpQsmW3OCQXg8KgJykmg0YIlYT2JWInBpFXZ0ovNW9ReH9ei1d95+xfY9DZQNO1
fy4csbAExqxNU+U/FCUb2so23JhPs1vF3hGNQFJgpm7vxLE3zTolOxoZR/1dY2AnOMCsoi+bHkso
CeHRbpQpB9u/ft3nSjgKHbMJNkpilNeIIOLi+JBBWXKOje2ArSKyiI5y/678qelDcIYeZ6y58mLT
iw9P6pgZbGk3PT609duTo038fD4WB1/XW0pGD4qaunKglKiRAVtfPY9805DOGP43otjrVIViXr+I
tQDcQKxAdBFKkQhtwuHJ1pSFJAYaIrt6IuX2mNAh/LSnR0VCtTaXUWMDsfQeYhMdsFpFHc4UPOWf
bvle8h9fZiq3Sq50i30Y7EqZYNQV+ENDUx9NXrcie65SXa8ri75gu7kHeXZ7QX3N3elymqiaVaoM
YMpJl/4SRhw1CsgzmYLS54znPdfHZtu4kCHN+NciCCN3C57KKDNZlUMy1Aa/mucI6e4IC7YISW9b
BdxN0IjkOdD/tMXdLpPDj5fU2Mn8TM4IVe/SoqdC8REk8ItEetqp+iLoktWhR/CM6qKCAE0x5USb
GuqA8ZNT/9KuT4/a8Uvy53lZQAN6FybCv49S2NahID8aeDtREsqlAZpDldkRQeT45l5daXKYpeSJ
8TRyvjonppUJDAXDqbMe5y6ksmB/C6smjglpKBjQVIbzuXeZEqa282aALTyY9GJqgPasMS+MlAF0
9GIZMgNDf05XzezNPzTsYaZ81KNGgc8PC3D7zOTzmXUwEQB5EqavYD79HL5oj8xX+EmTLnhHZbUJ
tlZEBDnVMgZ1ID9AiSHylwOXJmhv3uPsCer4wFKnTCRBrnLCJK7MjY4wmgiLrosHHoHi9Jg1rN/y
dS3TaddliG0vJfVdO/rmsNndWBXwYgdmLxTiC2dhihwnt6lA+wjQBMSqmPXhPH8o17rnVFKW4gDc
iW2uOKwPPjbNgdeRGfh7xK6ksJWkjixGGtvYkuN9ZHWodF6L3sXKiW+ltmddesJZygKts58izZxR
iFa/orCmj5p3WrRsnDMKFoyb67lTXQJzymlI3jb4QnI9tYgtK7YKAtMXzCPUZLjFN+DvR/BCsYwg
cGbFvxAb7U9ST8/a2LyJ3t3DGoViP+A1GzrGGsbJx1ChpP0aWsx9xVa1x2Hd1C/gkndqWGLwjjXL
jjhbcSuQL4YViBn4RkdjuUgr87asNChuUcpetsSZgnEAWamHk4qIjTbhvy5J8t6RlYmZPmF/tB3p
wvIRNKGZjuWaCEIeTc+jCMTW/c4vhDHqk45J8H6utaZecoooAyBEfe6m+Jh/aXZKMnpC/wfb9kOB
WraB7Tz2vbj2JyLDGJO1Xqe/7S9STbJmysHFWAcmSr5k7H5A+QpP5eipm2m68LvqeGvGwfofZzD6
zDlwx49I55TSEYgHTM+bKO1fvNlkLNw8tSpaJSXCZYgXePR7DaQ1nd/axIoGeCjNGP9DWkU/bfwq
YWspx+aakgzKqorx7msJ9FAk1NIGAUmRp1cgj/J5Q2aqHTS4pgEHnoYhoPvDKZtkpEGV6i9tMiQl
P48NV/vbaX4wq7gncrD9UA8MwE8u+fxS9nkEMZ5L7GHXd/3inEjECkI03qirFdnDtlHQpgW+xgvQ
qRginKnoVCQ73RPKtDEL2jlrqi+t2psE8je8r5tHF58CgiwVKn+VdH76WSq7hKb08jNZNgvD/DAy
QLevOTiqjOd1gAwQ9SIKpOLkgP4JZv/jW4NQ+YjC30yF3IKnIVLFVhI+bhW/0eT29Rou5kkFIAHb
zz8+kv4ui3imekCL/qFu
`protect end_protected
