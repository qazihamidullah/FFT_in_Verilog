-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OLmojF5jF0JREghDmAtqX1fubWzgY5hULn18HwLq7InZlcrNenUVpL67Jp/J6DLY0IGCzCUV8uBU
0LnUk5W7TNAE7WxoW0IBIx2FfaEGD4MC72rDat5f44LrZmN6phF6FZdZ7Oxa9B9QxkcB5qyOBCFV
g8IPxw9r5P/hVFhyIVL23D/vM1Uqsx6zRc5r51CJNF15d2bttPFgSjBxC/QsU0YojXs0g9vyAYMo
NcOSxo24kL2J1HQDa1dv1gIul8nXRZi4mqHzilq9J5croghoCzHqN+LWDNF7i4Z0bBtD1Q0aHpV5
8+rLYbUAd1PWU0gfek6C6tSfdP4I3Jlqqjht3Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1056)
`protect data_block
I+pliDh/U83RqADTlDuUS4xrn/FaIHTfC9DPZkL8fPlKLXiiUHv2jPn6dyE+KfS62GNPRTtoj1b/
y2i2DysR2nVpiV9i/58DA6e2ImhT9OyY3sDP56+/lZ4XiwnqzgkPzzaDhxyY/fGuFVR0K/T7lxJ9
GPj3Vu5NV7piVaJE81hQ8/N7lvD/xruY2GZZJ/iY2siBQipopzmLl9CVV7Q/IX972KKhslXsGz9U
6t1+yYjyuG6CkSX8lu8zOe9QDH8Q9TzZWACxt3JdFhylV76J2y6XYCyIe9bCQpMZf1//LUiRIF77
DH4AsuJpSnMNKxuhdnmdQXadGFthOZelJ0alQ91vpq7JcCciDZp36kQl/0pXsICTUN5dJ63FYSDO
pmbuBT3rdAPgOP5tfYj26288vuOmtxYJdAlY9LISRJsWLzZHfNA8fNjJbReQyLkLkUpNn3iAj5DR
3YcebpUTBzyjxTPb+LoeFteZCkiGdxvg6H9Ekg/ePPKdc5Bkms5iP7WcxayIax7rKaWrRL+Uhh2y
HiOk1RmDuj1IwTaIpybeSfhoSh50OGCclGfVM/1HXtn5KlSOq9GHm2+NMG9G7m3gRFcbcTo8yip+
mJx4boFkIgK3fjvIBqK5uAERUolnEPJ4/OorNzqZPz1GBgAy4pqmG+iBmPwi+Gzaymw5gPwMwxwj
XT9Frbz++N+Y6OLpd+LpdX9eM+2BacOWwMgthuqbTxrdEDbWbfWEjQHzZMf2Pr7ZWtcmfJEwT7RR
augZHtnvaKPUIyEM6RzYJlIbLsdS75rFCyVR73vwfbGXZJgIqujTwOD7zEE8QGHeeYwkl+kTOw+1
BkWRSm/BzV5Ee5ErXWuPSK1SHFPR19rbEa8GMxjxEXoHv+METpRKX8KrA4/S2UaaCiuzEJmEyoLA
ruPSk9LBz9K69QuJtQUg0XF+ZCR4PEZ5WtbJ2aeN4DU2YzuO0pjzi+L/yPcXtiRogoqNzlkXUlUU
GaPtm9RC6bry9PatSTQZSNIiYfOTZj/S/99PoKXnAG2wSAErCuSljT6GTjvcq19X/lGbTxkCLrtQ
vIgW97IoykN94sERQ5n9DgQvyCzRUZhlYX7KNOReWKbwgnRl0+jx2Besgj4w+riXhtAB1UHqzNhm
CNSa0j13eTjaAobwsGzL9eLkeNfXz+S6ZsWnDHWTFFAUMjAZyTzwQvmXH0O3PWHs55oK8VV9/uvW
0jf6yd/CNXiOMCqVlwN06fWhVQHEkJaAeJYTKKR2FuYjrQlWtdQ8XnUF4JIRz9Cz7EjYcRRQLGLE
scgT5odUVWoeQbMuhFhROaypNB9j5H0MN6j9kgS8fN6HI+3asg8lJe/DyeIoWD3eEzgqys3eUNpo
2Wes9kcFKWzQcfmAwrzOO0ZiL3LZ42ntyYjUfiTs
`protect end_protected
