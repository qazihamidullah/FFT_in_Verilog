// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 21.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
rWsfYV10RH0Fv0rPjWRKyA2uTCp+3Qr4kDKl6jfVBBdat1sirXCL3BavZtI28j8tS/GXpMcTpP2+
ZAOGPDtSv0su77cx4TvkvMaNvf0VM2nRcs6As88Hp+VtAqK2UmqSeL18kjIhtF5McBZKQNfz3Rv/
srs8vTq4ZBZIVhegKOBei3bBGfuzu7yFIyeqFog54LltOjDb2f90H94twm1NmrPTasvXlWH4CTBa
dbgDyJsYIHrm/UdltgV/Ma+fTsxcL815qOAYYzciWtQ36HfCQ9G82WbidCg89pbkS68UARt+K2v8
8XT5oa2U04M/e0F+xsO+tehXL/wECRN4C6yGBg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11120)
juYlAk/6dWeo5r2rc/lZqXQa/jScI7VpeE9qvQFu3v7uWNlvSnxIYIk00yy33EBpWNkvD0gPQRPn
CMuCjqGMNfnO/51xzOP5OC1Iy7zab8CRfPlDpE/wJzI+9s9VTuNdsCHhlbwzrFXkALbjfpYYwlHA
wj5Z6RVJ47kUJz+80OUdJYM7XQ82Up9B9m1TCP6SN4CHtjWazu5TcD2dlFtNn4lGQZTwBTgQs1LW
oGJfyTWK6vz0IxD63oz4I4U9Tbtw7aAGVg+HJTK6IXFoYn5nkyUcrC3dL2GS+qk1svxqH6TaDsiI
YlDny6m130iOCyZuXUp1hzW5OgfBesIp/8f2/bTPK55KQFIZlZ8Dg5hRAQLzd8IiYp+M5aU2ZFam
DhWypHykE52lMQDiO3I3tWVal0L9y6fOQuv9/oHuGf+HHxsho0UMHQ2tLkbCPiqv2KpJZw/+BGBu
uv3Xciariw41zjXZpN9ylvQGjJLTZtP/HslgcqLUYm/+nBC8EhhqZHcbSCBPfFZKwVp29cRiemCF
BtFQyijvvpojDyzV5kTTfnstYFo3gfIGLYCHK35nAe9LBbYTx7MnhIcuNMiGEBzv+tpIyNrhKWv0
9mICqzwzzUZ2MvBTjwmVki7TeWCbblJN9oXzePb8JbOISEDC2Q00ntqlmy9Iipfc4tddfqw//f0J
ZatqVAN6fP+UO/7jl2+c7qMk88udlnctghY+PuZ+qt+SWFxpOKtiacxPTLJJdug97/6dPm/1qycS
wTq2K/oew5GR22aByhQSeeDGc2ldyub+yyrDOYuvPRRjbCCtyD6eBJi/fRoZbjA8nir2cvlQr6O1
Lfe1eho6s//ejHh5GG4gVPvK6HlX5vZQwme4YAq5P5AMyiEpQzMO76QTW0e+XJ20h0aAlmNX6ap5
zp/14tWGuQQAU8Zy/tyjhDcxihmN+fnAptJZhlfWzq1Rk6p0KlY7qHv+DHdCoW0N7BsU/cvz+yJB
BfB6eUdK1fH57UsafrZk7VEbWuFufpd3lKaE57Eunr1NQTpVrDgvol3Kn7Ma2tY6Xo0VvNwn4cm+
mIQ/qT8eDHQeiAuguaf2xI8aru78oA66Z8MOYIWmtN2XfuSZEqw6JX+uLV0HJ52CkUChK4o/BRhu
gixu03dfveWEdfLV2db+syepG/XbW96jemWhwWB1kj+/C1o1aH4Dklq3L2T7gdw17rV5tP+3z4qM
Dk1LDV1FNwXgkUje726J4eS4SWg488ZDVm97yU+xA5k9L68LSrua+8hlyBHssYSCh4Xmw5RBeH/n
PR8L6HzAO+8lkRhapSMS1E2iJF8LqZCdfvy7PbibjDof9vQ8F8uN0v1Ke+871vv3QlSkXr8TeS7L
l/v2urfloEGSHydd6OzaNO4bAC/ljm1DdAFzJWjg+nkDhYhrZt6BSZG0vRcCYCSbl/3aSIg4UNia
QjNe182QqmEThoCHwn9tf8bU1xbnlxX6T+9L0KwGOGnW44z1eLm0kjO4VnKLPD+NEnK414CORLd6
Hzgez255+jspXyIMuq3X3DsSRVptguZY/Qpmem5Ox87rQf3Z3rYR4FwYQ60b3nU5Y62hUHJowYO6
4VYfvVLIUEoRmcWqT2UnzVJmA7w2pi/ho2toWYxSNl/1R7gr3KUCzcV511if4ME+IREViLoYL1B2
QP/9bztY5zeBSzqykcoi6qOLqtMHBY+7SK9tpMGzZXIzD+QMC7jpqlRnZxehk7wNKXANWkkX6Cqo
dZIQJoP0kwR9cO3TtkVrHxFm/M5zt+qAg6HAjVtsuWhqAV6Mws+v+pxTD3paiJGqMKQxN5PO3quF
xKvzzb1451+YNSRE1cuSug2vXNFEjYniBPrs4WiJC0rTrUNoJHfM5lhPk8F3sZSENEN/A5V7cgfS
RawiUJpZnfVK19BjgP9a2R1ZnrpPKH1BAbPrwIB5UoeZmdMMnX0fZPlRtql6ytjf3b0S+YEAP4y/
bNCDEcmAL8EE+j3r4swqap7HF6+2vgjC4WWwB3EXV7CTI9WAidLl5Y3V8QfCVP/pYgWHn6KEqfmV
C3uUjRzUsOFHm+th5cDOkFD6XcfZC5RMLFsrwEJPFYoEEC/w9x4ZMLmNefaJFrUWPNiApicbEf7B
L71/NGW0hlTCqAL1CYixLANUGu/vQi/ChoCfE1FCbwB1s9iCdTUeny9eCZL9sdvFui2c0yIu2BIi
gDfUHIp89fVHwwsQTcGRLdL4tA8sRvTjbArZtyHYbAgXBym9WSPRgSjk7Su38B61bguvIBMW6YI7
IzIoZDxJ97lUx1DQXVWHgTDULdblPIT1KaXh3/gq7wmNfhU7UtIJHJArqechAVt4k5EH0LXC7Z3y
kJDtSVkkwcMUSy2ibPya+h3hDby28I4xvNFte/dj/P6zvl79NjDakW80LiRG96elrewrk98HGTDI
+B9eYoa2vgh2LSe4fydIFqRk/fK92POpm0umlTPc7ENHswK0NZnRwy2+ujxO/VfrCYKoqNxE2hb8
gG+hW02lauyI5WIMGQXKNmwA0jmSMW271ATTWNU8fVJ3SLVIxqojDM/CvIZWgc8W/0UVV74tLoDh
j4t3bYn1HyWOIXPLTVwlFJa2Mc7C56MFBqtLaARh5/xxh6UjCMDyFvTIz4wfM0T9UhuBtYPvU5+T
b/EYUnTtnRzI936rDiVvZyliArpuM/KosOJ46g2+2WO9RfG319wX9+tzLWHMATLmogrkBNwD6J9O
h47f0HbILFIevhF6pcEEVQR2grOy4hlsBPXlw0TFSwwwlAQeYS73xwrnbhY1Po/qJt7CWw4zdC71
x6JdiBC0HlGA+mkfLVmNIXNQaDNzIxJg8eL10s1hxsF5Ukqu4cE4ZMXJrLBJ+a0cbgSn2f0TdYnb
i7FAvyHokCDoOwmjAaVlUnVjZAqJkpHQnD2plH5I69qsspnLqzfnnmhYMOiegdae0pzgNgHENwly
w01LGjptER14h+ygOV1wy28gzTP6BBfmsbikc/1bD6dRH+MUbRL9IuLodFrV+24dTygaXCCz2Z2o
a0u8EpTCV89UW0nivYHzjjy63WpQ0QFs+l3fyUw6BBifKlamXgqq6LWAr4BhQ4L+7jvAo3ab+NU5
+pyhjyabTezds++wK73zQgcs3cZESonJ00i/6+Nez4OlwuYgtN35PuhCUTW5if9k060H5SFOkgxh
jHzWCfjvMWpi8Z08ulZUEl+RiWoUL6N6uNudwuVEROqKWBZkS0MV8gjfjGkL3fkrmCx4OCNQEii9
wzjLevsXIBHyI69UV2OnEvHWXuF90+FtBWmWJbgacIwnig+k2fJuDbheBQisRueI/RAijYP0V3gU
a7AQ/iIhrKVK6EBDBvm/gvb3wDoe98ezZ0aXwfUnoSAlphlu4v+8vpe7KTdfk1PryQkhu+cFyDjs
myoAzXs8slz0eExg409CvBsc5L4YIVkNHZp/7+Glcc0ReWof/xpndDS6aHZG5q4GBtT48XeiKpxc
BcClBwIL6cRYefj98cQykbUPyRjTg6rfOzriAT8io8+udsFL3VcuwwJudMl5TQUvECnFiQzkvezw
hSVMApEbZ2ZjkkzF8iNuscCAbrYoEqMmvivULlStgNVCl9tHv31sM/WJs7HW2PdVOsgIFo3s8yNK
ch57DI3rISpcC+sOAZTUr4+gHuAYXyUBgmweCbvOe7ULEf3NwXjfanp8bbgl3tmpcwaC+bmp15QX
R4RK0Pg3wCkyzpI8OE7L1f383MaeqAy8dq2e8YbfLH7HHHc/TUtXsnjy90raTzqmGoDmj/AjIwcL
HVwcZcN4QMVfEzffVcLD4fri7TlOYZ2rb3MhLx5+E63PGMAN+opHyypUc99Wui8HX5qbtrRUPDtx
w23fPnCJKS1W3+lMMlC/QyHmQwfQ0LQSa2yQZLI4fEJS2Jn5LyMs4MyTOAln352MtBjQIZCrqDZC
yrpy2mSNVODRI4oEMawRBabrgamPzv03pMEaYgV5fLeMLPs3vChDq49IE1cHjXZ4KOdWle53lBUn
wwLX4gGi2qeGg8HwjHGaPl8+oT6BZAZDbmkk6gyg0VRvC6pu/O8Vw78SrkJI7UxVUy6QoSNaigMf
BBYQG9MOkx2OKMqR5SP5MKsDRdOMdIahvlops5Lj+Yp553MosncUzVqGS4OzLSifrynJ9mQeanr/
/+6fh7GtaPpOnx46mBOR5KdrJIQfg+Pp9tG4qUPDscr2JMOT39t6g7xU+eP9+PGXB61a94Mxw39l
7EZbnISySwG5Uw1hL08OLJEobVE13k0je8iwq2hFNVu93rXyWDFSFvyKPyFErImdLi3uwD+pCEO+
uWmYycr+fwG997L50vgK3bUdosQKE8ug5cdNff7vU1l+cXMYM5CaZgH1rlJjmn+GI+Sdo0UIVnpR
Lkct+52G8PZdObTaNaTa96d3NK8PMMzP1U+pcIr+jETYOCa/+jA/S+GVQ4VY/w5XFwIJVv2CkVqK
bI9oL5Lbae3mcAJjObf3b0LN6v6PorevgjkD7gYvuVEyhbhgQYYW6oGcg2/nkoI7kV79ncAho43W
p9aqxXBcmeLQrc8Y9a7i3mhykBIOkWp/xAdF+Yb4sUyFi/pnu0tIS1aFuYFsyrpKyWqtfOzI7CGC
FuDgvZjS98a83uL5u7wanptGvIapNep65myeFVv5QocPqRfVfzyUZEGCUc7nkr3sDaBlsZwwrJ2Z
+gUZPj1H0jHSYPPIcRDs1vfEI75QSFltoJWYDduRtpVGOot1abvJcc7NprF2fzZq46mXEMulvQrG
/9Zxc0gCy5ZRVBha9h9TCP3qFO19of9989v1KAy/H+K7Pp4G1B3Ls/1w5GNyixlrgg0OcZEvT2rY
eXYOwc9qTTeprd42i6US1fp6e5ixkKNYChULDBLziYHBP/SYdzJmR3mLPjM/hFLVKZD5Qb9GZuFu
FoMy7vB8HFpY2tlHnxOB8Q/kJfx5dpjbCgUEqsLPge2QfkBIaw9y7CTRB7U5JCZ6CZaBgUzvxK4I
kqteFXGqltg7OzCtBf4P7MHitqatZ86pqlTR/p1uWYNIZra8HwDgGpgfM88HMzcdOKz/7Xho7o8p
NFUjlNyP9VH42JjkejGrQ65YvWLi6d5PUiQnIXlX3sbGH+ZxBRXBMGwyg1bDoOU2zkfm/v5Rj/Eh
VujeAsed5mlFm+FTI3XSMwTGsstT023dVtqWBPnVL7Y0VjhXXsCGJpkEf3q98AQ9uweSr4wJJAwI
4gIKc82kF/NL2lRUtTOsoG9PHNju0rb/9BeovRY9NTff3i8O/eotmY7KDMo7QDsrUUdy60Qw5i3+
xqNL/A6Jxh9+03IvtupUpX1UROv50belSCZbJS0L3K9hFFYfPZbVnCNhm+GNYq8xfyCqv/Xy963R
hjPnsjmibu15IVzmCjvrwszWAcY6Wk9s+b/Dwzd8cctaRuqL03cE9kgTNCq2sYG8/GP+e9kBBTDq
BjwM/P05Na1nnAy+rme6BTvGbmlhFrfc9Sk0hjRH7dMLutz4QbvgXZv5bKzzFk+XE7YpMuvYzV8F
c7unE2mu4nvWuSRrn8pe2YPmBYjz4m730NW0fY7e7bkPjd/+XNptYnc8LC5Wa0L/F89R7/J+Vpze
6goFx0r7qE0y9nbNBOJSpKaht/eee43EEFHIeeE5/74okHBiRTOFz+qrISEBHGQ55DdPywSxxeBi
a3axOFTw4eFAySNSd/1SHQTUYLLT3XQ4qcGmi/6bhEip3B84fcgJHTZ5zymdQrtbllshrV3cXg1H
8LF3xXEjcGbeL51jvrb4HZZyxdEIjPZ622Sz5uETaP2fum0Q893NzJR6k9yGJnsk/L1oLwtAjD8j
iVt25THldtksBdZ/0IAa2xA24CvRa+Cof+oV5693xBy4MCTP17LGilIEfi45c9AxLjmj9PbkfCjx
5FzeJatK/YII0ZuYz6yLsol1aWCfoNqMvRfM0vPB3o6LI3TIuGNmIDT+3emQTvFlqnOffEfovIjc
JPCDkNPgArHGxv+lMiZ4cri43KRNAfyrevvwHjviL58TDfiNf00+fpFBh6BQRC1Qy3rZITEawD3+
nLNmI5M5Fq7BeiriO6YBh0/03Z6QhlETDJKNNqWHG7C4zgL+85tfsHchLTSgmFsqWk7OakWeKkAq
51pFhDuTOkhsXwc9h7n7B97yRTBaAWsN9MZokJPZdF9br4Xx6z5PS1i0WqfG6tTCJ+XMd9BRjs7N
ifAHCCHiBcpggiN3UIjDgq6h1yzEtCyJXxZ4PrdzFdg7qyYUSQGKNeHr7H3Nqwz6NwdPdRUl5/Ui
ZhAyC45z/3STRxrouFf6T10MnwMXrMipczCXnNuV8VBZKugo6txdmAqN+m2xXwv7qDgFgsxtrc+D
S89ejgbITTxYwbasiZB57B5Dzr0Qcapx0MOjuXlZ721Auuc9xmUQ7hoFHQdeSTs9TwT0hD4a4745
MLfwkC2YZgAs4smmTy/1mxZfJyBExTiIyr9+/yt4/zMVyT+cSHHmf8F/4PE6hCa/+VHmDUMUE3TU
H1v52vvywQFfmhKCyfr+nEo7w/pD1RCPbCnpkm0lF9RY1DhZLzGla5c7kdofX7Lb970OZWF2GEju
7ISrKvjJyyPLMD6FZtQsROfRVrDGpmc1ZUwbObQyDDv1Cv1Myx1d8M6DcqwsR2MouziABG5IucJ+
tOEH/mar3iz/JmniFqqe9qO5S1Jr0nynztNTCPjHaYxVugoO/fNQG8QQKA0YreMJxIAjcfpuf+7c
7ArTCBCvk44dXaUuFOKYMQvGTE6izYU8jxRA7tjwiKPdqS1flVQk2HtogAmifBQdlu6PlmJGWpwV
LbnJvhnuUf9uS0u5zoSnWmMPGOK09/goM0Pzs1IoMH4af2WV+T/W+rsbgdA5lpWWm/XZGvvj0QPW
PBAjctzmDLrFnSqOOZBsbH2dYvv37LTBOFO542mvNhaGxZDzypCXVJmkmVngUvtDhH8/a2tfm76K
LTr3VRIPRCbN3wqmset1Y8Ufv+hxq9uPo5MHt5n10XGnTlthUcl6YQliC+HhoVv2sroIU/l7KZSL
FO7xIJLHbbmMmGIWbtzSCgqRz6geDo9Wpewrj/UYY5OoFrF9FTICdGT+5IgdGxJqsYgbnSdLnwZs
LGthMtgFoovuJ6ONVxJYqY+xwBcMPa9XGO+flvyNrgpCdVP4hGniIlpV/08nuCxIkRKJAPsDwgQX
6Rvpo/coZg41FlrCCnW4Hms054nghlmOshi0EgU6u6sAd7m8HyUf323/dzXtexUdTPT9YDdevAVg
VgxYv2DY10MtxP2lBcrvXuPZKxrwJu4HoqfBzcfQIBkVXYiYRcPl2FQNJOA0TlsXc/Fgs387YoM4
JiI0JC6R0kPYamCnsJRRoKAwsLRi+jRvjLBdo6hTX7P5S+DqPApXqv8Ec8Kb9Dw/8V07mRAahcw0
r7lfflZhFzyjcyZFHK91UZjP2JOwYMl+D5bdt0rDEPIfaiu/6l6JYxcV3pzW6J4KrF8FhZmGTP4v
qf6eQsm40l+c7iEynyU7dY5gR276fDXT7QBvTqoiPpHu9vqJysRs75tdfOlX22ynBdqzWaKF8db0
vXY8RGatAcO2UcMNNrj7Mx0MxRxiyuO+tqudQZIGj2WLXSUr9wvgIHTMmCzJTEiC3qMB0OYyW4xJ
FnZ/pG6LoXRKF2Qp1Jpd+zCKqLcxAcUZpYKkw07RxYeD+Uj8Ho1IHFnU4qhTSvNh0gU+Q7WsN9cj
VHboZtWXMtEnDQp5Tk5xpyshjEdctYOIVVTPwpFLxv3o5rm4IMruFbtPhGvNGtE4y/iEEggZch/W
F/6eKwoud3b4MO17nzqrpJ0s7pb94YNsnhN9Z8rbRWsOcRAG2ANKmcrs/IknVTKMiB2BvbSSCTxn
vSChloLyDN9UECYC0b0a57NIBS4Yt2hT9CYseRGhGJQZAdCYtsq4Hjy1sl1uUXknY9Ds335bt0sO
TNZ/qKV/pE8wYjl+qCuz2Nt7kmbu98VautyEwzT/oyfNue/Lekw+s32kNZ8zSMrXiW8hTvER4B5V
Ls3VeTYUKImRpNiFgaGayhEs8XG5TwO6Jsv811dLvvZQbPP2eYfEr/FlmqZIVY2T9u4r34rYEykq
YMq39iyY+bZVRkfAv2PCOCGoKGwmTOmED7R6puVqsvQsWqfJvuX9/om2/5RvOKkG/TtZiR4N3n+h
pNbctWKhq9NPtmhSRYnktiZw9rRkVHysqf/MiQ0UyQTEVd9S2YLne7PdCeAdUvYU2uytkoKfUB49
xFjj+PFhVfwoijHiHvToVngAWbADhd0C6/3DYbbIQYw8CevjkPDFFBITsZUq94OfOiyZBvqOGWb3
+zj6dUT51BCAy+SeLQ12yfOrcLT20d/YHAWrbQAgDp3SoPhyurWdWWAHrWG8aPrYTwUjJKprqtqk
vzOgYZPvjufL9xw4QOA4EZ4t/MFr8w+gq6tQqHsQ+d90+dBMYBPQgwDMV0BuM5Zj0Bvi1fGZoDNg
IcmNZL94Szg/DsI+VRcePc4kNc/od3MsJVYFKeiwJcjSGOXlDAIVqcozkHEfPsrg9rF86pWm1dMM
f6Gc25KRYySPBXye6V3wXQzHkBl2KMQ8cvPVOSpwceQoxiKTD5tPRWlDuZgBK5AsgbJXz5bOb6SJ
rs0NcbaD1V8PxMffIuKEyNG1ofKyDWARntsFEtnZ6hNkQLLBWSlW0Ngf4NJYMojpNeBcsexTwK2t
zefBYpsStD9DEYSCPlqaJ2m7H/wgMU9rriT9x26MURbAFzwq6MckvrzwOtq3rbHPOj68140SYO6D
TyknHRRDl6ZT7nbwuHqoSlgXbGKsBgQloZJZN79mLIl4Cg9GkAa0wwDUpTB3aD7yr8VNXQioGemg
a3c9YkKnV8Rjxz++sWOzfK/ww2MKF/4JqayN4ZYaYj1bgpIxL7coH4N/7vZIXbweuBBjVnCAQDbz
mCdmM+OmN4L5GbZIBXaQDN39w2t7V/eDTWoeZeXAPkqzSEdd3UTaKjhG35oRTvKkUGIm8zNhmFNy
kkB1s2SczIbm/yd7uEXpma0nDt/VeAIcqBeSQwculH/Sjzyj7RAPad78MB5gHp5B+6BPgO/Tw4Mn
hQLME5RWDeUoCbeAUvMH1wGj8yK9pPkxhQ5G4CHFLXXLRbOCcKqki0DlRvnJHmKJEcDL0WUON71P
y8tCeG//yO9xzIYu/ZWADoiJT4y3NCYIw+eN5WLyrI/D0ZdzxQHHLp1Y4DnrN8haEASErLoolif+
nN4NE8Cg8nw8ZVmVytR8xSwN0EPJI/KoNb6GsIwrMrzEKDZV28UKicrHauJJkuCFtQwpVwvhaJT6
3dPcURISm/ocB5Vb9OBiCWTxnqx+s2FXlMHj15mM5T84gk52JG4ttVbkM+eTXVkH9LRU7zZSz95o
xVVsexOM8OFrXmIYuFSac7L/6iTrFhkGcbl2f4Rt4+jkHxbBmmxR0VoHYFGwRh1rXQXZTp4GLeZ7
YTcf4RG+hflpXxUgB4qgaRIeF/IPUnPqOj0goatuZdp8G+fo8UhB4A3kBf/+tQgxM1vYdypnCo32
v808Du+OBVxm0vtnkKd7N7651YAb3Niq7A/zwjspMKUTLRuszhn11rSrCGeLpbMdnuJcsiVlkCt+
dTM3XFVWf7xvmioEpz+yn6CtkY2onn52c8ZZiFQiREq4YO2lBpQdEJHlwjbBI5nfbwFbn4ukuLpp
oFYnbTwiSOvti/jxPhU2Xfpy/QgPPhFSXV+o2LtJlqSnTD0DrUET2Im9wdLMe8UGK5p5thRLKyfc
V3AbDvvYe/DF7W6jqgUpOyjNCaG1ZviDJz416nvBVlIlp+wZ1zvBXO1z3lNQaUG7JOPjceId8l/P
WCrhLEvJEIdmfc7IQn2vfj/HdZqxNT0B0AeCpuiQx/RDbtE/0pfSRks782A6q8eEvOFVJdo8uOIr
D54gqS/p86nT0iwnPG/hdJ6yirgSAE+tZv1eYwamVQXI4acX+UOVElC4hvUr1SbAq125oSO4YRx5
N+u7QPwwvxQ23jd8U7oA2oOJBeCvGJS+kp8frhMgusRqJF4NcMl4b133BamT0Eu4UlGsab9+Mwc0
UUCo6XtOa3qQu4+ZfFH+0vAsw0KhjEIYZxhV9pXN3V5Z0AVzl8Z6hdYuyu3gBGqwbOBoo4VyHyXU
kNAPtXoaXF/93gcX2kFWCNEHO4AY3pMBUb+6wfhEZ2X3PfQwby49gN6KtRe1gA5WnH8eEGv3AKON
Mt9W1xflxRDCOS6DxfpJKXH++g9hEfwcdTr+iqB3H00jMBupBROFJE5xnrtcIYfRBBHr3haI0RXD
BlVH5b59XXLij0XwS3zHtRniJiT12fHb3C+DK+0LydUYL+qDFmeXqBb9r2+6AlB9nXQrw62cnNrM
KqiwRQu5MmfWEYWpadBEJGcwHkAz8JqOPVczA/yCuHaMahk0AzEFHkGu/3gC6z9CqRXAjyFkxAhy
sWUd2vGnqkKTFJ5n5E25h5C9nt3w6itAlr7ud11BO5tx7mCwb2UaEi9lQZAwBf9ak0SO8rodDvcN
JdJgLtoPDUgb30YzH+0iDN1e/URHxsmuXLbtQqPQvNV/N+WbX+S7uA1IhEyuHlNEJYreLKDP43VR
B49ELhIo4yE7SmS0TbhSbBdte5EqLm/rewBjqMhfgv2txvW74ACqMX1NfX6R0J2V8S1z2g9/XGfm
FcPIytCuIeEM/X3zotB6BubmIvi4GMt9eMwRKYmWHQeC1G0jqe4XbQxZHeHb0WpSXmZ/RH8Gu4kg
FQuVr0XvYwc6HYXE0rE0D7R3Pr8Z123SNRC0bfAIGXQS9ismdHeujmmjtrdJcqDXdfCKXwg5h+jJ
K9oYmWcRiJ7dj+bp1c+0B+MvjWHrTauvXRADOea+MizIUz7+tvgfYuANPRn/Fl1IlmJD1yDHZwn1
aXrXWtzoQRblw4AbN48/Rkk+IxcCx5K5JgZrCBNapG1KOcQswKErseRVox5zZD9uObaNu7P7Clci
UrdK7u01Fxfv7ZGpZQpzeUyIQL0khZGgU0EinQbp48Z1ME8ESy8FzUPCvCX8+cVzmrWA04PJqyz3
jOtPjAKZgKStLw+cvuy8C+P6JO2wVWV4eEwHkiaeoHOOYU6/fZNAs6dENl0PnRGHdFI3+uemaeSv
pfhG9WKe9tIRvcshc6Y3VjPyEnGWHqcThI+QuOgTb9J3O3jwFxQcq2sT+C1xXHM1451vMyYYXQGG
0CHPF0cFYDGXqQpxPXbom2R65fA9aoYqShiPjwB27k+yGyj58Q7ddA6lu5iJt+rXKkk24JfLUlnD
rJ0fQilMum/3SdHSYuCt8fTGN3AzI68SpeJcLDViT/hKFvR/44wjIzUZ0EsohXW4c55jbq6Kckoa
i8gHyWxlWs+tKr6ehKyfL6sEPJczopCcMYm9yvTUH8H6L1d45WeDuay/LuhQUZCQtWZpnItdvTLe
kFYa7DEcwB/ALLVu16zrbh9CyegGvEBKnmKBknLdYup/wAqAzhnsx1jb4A4HMuaKGVp8AYJ4Iz+7
bILtORu1DVpSIQvhNWm10LS4hXldnHrkhrKFFlzc8PEofyxRlXaIEmgf+zLz4BNan5p6aUVxbYcN
S1IKO8sfHvA7fk31X3o97HHuOLr4/FTbcMGe/ZY1aE4zYo38xufjCEUTN4/SW6nYcrxxAMGHqLjS
gjaaHrgRhXGgBmLqYxACqWuHRgSZX3OFp6MJEyNlmtmenosWGwDuM17f+rjpe8/qaWv/QXU4dF1g
WimgTqoUyKGOH9vf1MEO+oVZJWIZrI4S0yHczAIbTVJqqWDfG2XaAezGfKLA6RqOMv0wa/DErzq5
uBPHQ490ZjsSEent/O7gb52iWv41r+O5c6ipJVLuF54IW7epThG0oG4AhUJUE1BzgVS7kNWRta0A
KD2u91jOD1pT64wLGjAooDoIg1aqzICiCQPwynmAG1kMku02mkiDNk7DxcHPLoqiuATZHUKv+yUM
owYLlzSJBCz8Zwl/BDfNoQ6QFoGbZIiWA2KpKk0uT0SMh1bH6kTv5IKjJpAdYIFkjASCGKHT2ZVb
+5fvT98+x5Nd8pQARqW06aKF1ypI/TX4pQgg8zPWJlcVuEJOnA5ugHzAdCzD49iqW9y20A7+wrqL
yq6UxEptEnHz6ySwAhQwNDSgfd0J+Gaz8q6psXGknqQkR9RE0r9DZPtYgkjM2Ik0TUouVBlE70DT
+0l3g0uNZS8heFcLaY4XBKietgvZiqFoAYDDIyaH/QxFi3rh5ulxKYK2blb3YuZi4c0g0HsmvhM2
1tD1j5+Vxq3GDa6jUAyj1aB46wF1jlMb49U0yU0+wdMnB/GD6uENRgnvq2qUVt5Q5ltwaOy5uoDC
ruQC7Jh99T2rpQTyQMBCu08AAYTt2OhD2P3IpMOJUDNoemZin3BhROh8biB1cT4DT96Ou8pRk/bc
hlkC6hTV3InDmAhnC/XtRWBu31Z7dWjOr3XQcFB14WuF809EVkjd1aIp46NFbztuzTdTJQRDSJ57
9Wsrxn2fzKTuxwbOnfkLc3gD2dEISNSDTI6yhKuFTt+APgGVwqAV15tsDim2aYGQO0Y8WQk8r/Ur
qF6/kA6P4GpjCXWK7BFzRMEtXPnuCWy3aDbr1BNl8TkvUSglaMkPL9iJ30QKh3rx/HahIV4ePxd8
66JfIGLTTeqW2VLaz2/2dMWbV1iHsZ9Tds9RLg2H+0pxmV44Oogta05pi0hsNanjBRdt+Ipzighv
c4UYtgbX6eqRM0a6txysQYu1rHzIeeOhnYtyHK7VlTtSHwy9g386xOiQVve9bNcMQIaLR7CCTAZl
AbPQvnBCpm7u/gL45zyPWjDTdmVPT3meiWCD59V7gsFW8gfSyIjNBt1bZDjGBCEaDzlgLmUTPBKH
Rp20bvjCuu+z6JFwQwJE4LPpRk6YRj+hHexrUd+Qy3rlr3jWag/cqWv+bo19Tb/UIW+WAfAfH9sj
HAdiapbkb2hVmC9W/QZ2sZ6xyRaBgc7Rp7ykg1P67VdWQV8ODboB+/26zEyBz5rK5Fe5qxBD7vjY
sAmGVbmIwevWycH4dl44KfkDTJKpMel6aysY9IgTdeOmiFVo0F77l4v0O1LzmU9TGyBY96dyqxZa
o61/+qUYPr4Xlrj8klD74Sk1mmI4JKI5yCn34mH/ygXslI/rDACTwQTOtwBLhz27hHrGtza0enJr
3dwv2ZHJm1ee4A1bed8Kl+IBoWeJsKRm+d4Nd4CG700Cb4i/l2izIuP2o6kYXijr60PRHcfcWmzm
1pTQ7Rizmp4WuCBSi8gzXVWLurxQoAqauihNl0GqxYqImBjKkVB3fybIhgv6ZhNs/5rUtaUGiG5T
1+K3BRoyepBYFrIteRJiXo/QpKDieO5vPZVSF/Xs5vWWCmY55Kb42QfjdfhTEDG/9hW5YJAud7sI
qB6QX1mYY35ZtA8/6kpZQZry3xcnqcWmmaKfmBh/rcbOc6RWPyuD76kuDZ8fK6PE/HvvuSwlcBcI
l84a3uIMyZokA2uzpQLsMuGy9AyVOcVLnhU1yivWYUHnhPNEbA8GunZ68C07Zvbc0X5aEucRdjzO
b3yYfyAPAj+TmVH6g7nMXzd/umJNS9eia06W05XRA0ha6vSaqKjesMW4fF3P4d0h+5caKOFUXqNj
FgdQ9GVbyeeQcizqqCJ6ldAeUYWecFQVVmEN/tqYgusFiTWZR9ZzNSpmKQWtd6k/dgFkTUCKrrhD
Dp3lTSEdNRBEIHm1AjyYbsAQ/BkC6iIxbdNjsj2NEu1BOOaWkLaa4PUTiCYPNoP1OBQAxag5r+nq
psJaO74Dn4ZQb9da2RbMh2CrLPZkQdk596s5mwBjMEZ351BxyKK3hIGmofV3xTqsdAkeTanOVem9
b2BcA3DHwZL3DcJp3j+2HTFIzgimErdowUR15jx8aln2ngZ5eL60WlugJa8zLCh8d8atMlUbXNEi
lC5mwOQTXrOvNXc2BC+hVPQlVnD5lL6i2e5GDktj8ibZxb0XEqiBdqRr5NzR9zKMxPWDrk/NixjZ
okEUAKqvaThEFSQg92qpJCj4GF1W4MHb5gCcPDwwI24FH4InCrDR1AO4aUJ7iEgsA1AMypQJJy9K
tnHpkkzj/Q+98shkZKGv+2TWDm3yv3NVCS6XoOBxyqFP9mK4XFBzAWltdWavHrEMEdNjwm2LXIXP
OyCaMzjKdOXlBwjl8I5OWYP4iZLTMGLpjpYEHBVlssvPfiWmJ90jbf/+Wiu0SG8W+uJq47/rDReV
RUYaXmGa4MiLHKOUxS9Eswfnijqvcrdi8JtmnfH5FcOzJIFhGG416hBj2LjCtkwLhE6L+ZSLAhVi
Jks8tT1jWZ8arv0jEVqeD1I9MjDE2Wc87jYuG/umhg1t6yPNu4Xpbh5GIOZgSzx4rkeD3Hu/wo77
jkRQtkhTWVXnxQsu+WI0opcgv8b7FNLaCP0TOwvO1xagwsoDnids03SXzPU2EgBLeP56bHpyeh1Y
9mygOWxwMZftH+Zx5/9kPM7/z6b2+CXemXgiezc/KcG3ZWBjrys9lkJXI9L39aEV/56rGmscnXKJ
fhg/9aFgBNRfMRKwVaMDZpOw05VpJYvcMCW5LuN2d6G/8kc7k8w2ipPGvhsIfuKklFT4fjZ7FD+t
BkPBToLD3UjXRWj8XB8G3I2bpNJrk4TlbRUOwJZVfXCaC1ccd7vMQ3pwN++5iohc+7FtXfRFulNJ
VY1Edg997YW6H7VUEhbDNYJQQqZ/WnK9YjbPV8NpWR7l94CxPPrebrBV6ibqBpEkc4G/HzPGsE3W
dDAnogc=
`pragma protect end_protected
