-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
15gSppGd/6IHkMzo42kYCLhXAFgR+MoK3beQCKeGYbeHebxU1kY9O3WkFRem3TkvSy5WdfB0Ckyq
goON6A2fraBI7Z1SkLgNc7GxdOaKSSEeRkCnOYXgSJJSuAYBNuIyXKkk6Ezsa/Rzzhq5F2xaADpn
pcQXUvYzMLZJQfK1uO3mZWxgzzwGzvOkz0ppNP3mi4DaD/MaGU+Nj/y3KbrYbA4PvTJS/HMYvXY8
rRep2TZRrfWvb5vf6sLb48FSCgTUV6Fe9OuR6SKPXyaFo5fNMD+23xwLBRLhaz5i7M5le9SHJu01
E9MkKrJrFIHqXzDZ1+XgMZv+KFHlHEIUC8Afpg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
OL3Q8YiPlobIOb0KRCZGRKyVYqz5FToiusy/ALY4KL0eeUUhf5LTRXKjK/4G2exubNndYcuNp5sv
K3a/8iYRfM/1hOxUijCt3dChwjCisK8Jdqm69Q5HESZMcw5razsE8zZXAcKmb64+eDz2qbi3b9K6
6sVDdWS8JD7gJlofBDXaZl40dAZ9jNhtXRU2Ad8FgDrfCJGJ/NdFG5dBYR4nzTCIL+oJGUZIxBOi
67CMpAWQiLj1pyQLtyxeJbGmpmKhfb21RmUaNbZ0aomFGzKqjDXMGyDfXrhvRJuMbs2Oq/ItVoXN
ZMWt/dym2r2i2G76vNoQhVdBFcDRvr2ba8dB0RfSR2db+HnD/iYqc0HaWMXxiLRFYHXPVp3TASnw
j0IZ54F0LHZDDTJzRxLhu2t72HIduj4J3z5JeUqjOovuhSVAF6SkG36N74a+77SIJF4wY5pLFQdI
p1Tj+xNZCnJqxQGzVViEnJI9MQzZhgGAO2Yu3Dba9xaYyv96RdAHa0qq44lGWaTN7JWOTv6jaUY9
oF7RRtPKksL9LvR/+0QgkRBc+F4wgsqOBekXEdS5EzkSLnpXeyriyeoxpH3gHUl78PLH9gq1uG6Y
+V2RUuFLg/tet3jT8Tp01tUmcqWWItGgcjXJFZ+1sMki7hN9WTw/JAARxs4g+QY9esSYk6r3Fu2S
EVIFFJ0Vs0SCfoJ2pckphtPnEdREXJYGPUyNKOpNAzwuUXa/s5QhXcgy8bH25nrzwLrJDKC6RFfv
F2O+x8HYdF/iuHIjCi/00o1b9a96aUOoTUXn3maVJg16fxRJJDpmAJT7ltPcd0FqazQ8mTft57h9
sBvxxCtryUYQFPALSEfcEL9m07MSw1Wv98RhgeurWJ2CuAnA2BZEhBCxGRarYS7Wymc7Ar70ut2K
jiDAXF3D8/FFatoPrqVh/ae9vGdD+1Stvu6bjv8A9/asVySusCkbJVkyFrPuRoGvDepGoHFK+em2
zWkojx4QlJkh/9pOGARLiWlyUIvK8BarfHkL25cgbctiNyv7kBmEkVIHXWv03gCrGjjRmkPCIwY2
B3d2wbMagYVfJDI1xZtu36w04LxWT+pSswTnadfTw5IvLfDNCx9irV9rtcvsonxdHcMWuvmpaCwF
evrcKgdFQY2Mohrgkbl0SIIeroSNtoJf+FfBVaZbNDzpTlyf6rN9r2ujdsnSg4XPwd8QhzgfJClt
TleipdNQFEgJhd73coOXeomL/J+ju/lZZUUfI7PqIRVgxRXQsDDWjtTYKyeGZKjbxA0zHED8yRO6
QFZdZlQQXQUnlLfuS+6f/n7S5P9nbmNUlHBxTjFtbpQa2vvLeZQ7gN2hM2cUdMfZhnfUAsFk62/D
1BazMRZGCuaiRiLOdNgqABDtPxw8xlTuJ7leECbE9r+lvRrZe0isvFmmUwv96o6pmKrfbNa/Sp46
of/I44RV1qYqKcvqRSN88mczrE4Afg+G+N616Mwrk8Zfx3coPPAakegAUpXZrKM8iwfl24oYt7jc
jHO/HTwOOAVCqsR9bQafSpDaN7VHz5eEqfyJd6uX6gM7EMkqmfIbVXCfAtJiCksf5BsaCxf+X534
lasM9FdiBBl88w4r9cM7PWoMiHKae8xTv6lAKc4w8QZe7ts8T2PF20a5fFNYePLfmgS9i6hWUZ+e
V1qdTxJ+VKpcWULQ2DtagbsUyquRVCP2vdFtM1vgWUMiZ0mXDcGo1n8gmRqzFWvvOpcyyZ9OIh3M
pqm6FPpVw2DAsN2gACYdvWBNg30Qp/1mDl4fG4hdmYWTpi8TBn/n3MGnVIaI2n+hWHNrwbiiO9u8
XLJOrZsTkXDQXZOz9zRhkTj2U6R+8msre0lQtozcPFPjt6aDjZgEPAfoOMmsKL1MPoUgzW0kUT4i
ii4Xbp9+Hn5cnA55D9b27J8Zw3DrGZc4h+D1gfxMJ4aFv2LnBEWOgqLcJct17avV5TwqJKkLO8X6
j4wI7bXMm5/BVNxSEXX5bNQjc0eXdpDOV8xrkVaB2FMmLWR1V0JCa4HoOgVgIqzrr8x7KsgGnG9n
YgYzqrutuyCmhfBHZai2d/C+HIBBtTQDSqovcGn6ut3mFAqi9c7jejpjulHG0kHTZG6idlc/hbd0
IkEDptjk4Z9hnp9jZx3c559U4y9oy7/RsvmlvlQ+mBxGEl5kZ+REMimuYV8b2Oer24sIhz4u4kBe
tCQsrj2vpuMdN+6Loe/jXcdP2ng5BZpUHRFRsJir3LnICuqzyDNN+LTijSjLSVUxTELrVeKOqS/O
7QHB70GzgrB01/xli4oea7cxYTsYv4s1eoCG/6e19fECG5SXZiwRzHjoYZ0rGEL1HCLbQNeVOwO/
lGkQBLb0Y6/vQD+UkqGvAsmdqY55NWS9BrplYuKytZwCg42c4vb9LjBv4bLhrYNwe486Fjs8c4yR
A/vP3bwslOuJQsj/rjxZUskHlX5icrVqIZVlkM6Fy3Hb6X+Rcqs+Yo7ZH7NTL/RzCF4dnRoklTn9
qaHfxYP8d28qFgdUbQfqyB7Q2t/vl5MgynLeb3nDHlepFq1xuCnqSkzIJzs1CG5pfL57lrEYTNmC
hbfo0RlBDRZJ4iA6pnZ4Dj+SFY2MBNojUjoJmgcuTacezP+CPJUr+txeifn2PytouVjLQN/618BE
i63ij9/+jUFApjiz+TeO/3aKwgbYk9+/7X0Gw4zUOs5VpeHL4j7FpWV+R+gZgWIqcQWRY5D6XAv9
QMSOkmS+YFNyNMmhMs091zUNOoGBJKOCFHK/qwEwHPoV6kLfGm6kXYmVFgo1VSXKxOT+9/vSZDCd
YSMdJYM3hJarjhy2xdWov7qG+ZouepE9dbu4TnEldtHmB6pH13PLYZKZzYCSEBRUoaa1OJtQU2yp
tq6IBIPop6xKRs/mCsfmMW4Dmi2a5oSZZrE8HpgIZaWMlWTUp6BmYFz8FxWkpEb7F7i5jv1rUg6O
lxsxkElc/DBVgSGpTkVmH9kBAh3xRWVo+UzxHzxvRR9KMt1oc3bgi116AKmACH5ljn24vCjHOLR8
81OAwSWGbOy3C/7QGEXC+V3vovU013cC05ehwxwwYwK1KZPRDEqPvLIUwpVCWDZW+41JqtfxnUOe
S6a8/pjgnRoUmI8FmFLqoQJg4AjJeflsxlRKZMsemuesmq1slnSZPMTyfyvrFHPUCDXcX/I51CEM
GijZ9Ez56V9StMg05fCjH8Hei3wEHoGnfu6qSzBC7WtH1+s+KHfho6LVypDuT8GrwehzxO4palsM
UgPXtUuoqIG4E/VmW6cIk9LW4Vhh8ZUn8pwri2kchXAOW4ThlHwS+d+A/AHJhASd0fobgH80iiI5
aTY7HpTKUrrgQDuyWOfKSY6b44GLw3l8SNRpMngiOxsVl3EeDFflc0aQIHTiLtrMXivNKfbcLulF
f+VVH/xIfW2vZMOu68k1nF5vCA+PAF9D9Cj+unkiAuUR5+Vs2wDFm2PI0f1aB8vXNAvPf4MWKKTC
aI8BOheBHMoEnh6ERJ8MCy4xhvhpIXEEn9Zbcyq+RxKnbtZzzOdgaxTM+Mo0lvKLJuuFRTeQ3Rpv
lDjMhTpas+Tr/BMD8ceWOs6mz+j1wYRy19D2B0I7Ot76YhCyLmxxZ0pAS3cmyavrpc0OZsR0sKxD
wQyFp3zSKGK8oZd9j/hMX2WUtsvFS5curfGguwd+z6rVXvx/S9fi3Zz5W4G7pizGZ6cFahqJvy8u
O93R235/yt8gjz47gFl/HEC8mmHif+g3nzY1mXhMFyU87bXIuqkPnZVKJ3P5FtMfLPUV6xUGRJ4D
bODLE4z7pEYEU9bzV+E+U46MnClNi2N69afGRbO4QVDgJnnQFsC4iW2gSs4S23pFOeEAV16nIGNy
aLMUJpm14aRmC+CoSbE0AjGA+aiUdKopeKfI9t7bkdhHZkim/O7bYad7KWaXEl/Y6Uk+YiT4R4wd
xfkOneP1hN/cbdLL9mPHrX8BnfTmor/8cC5TBVyTZx7yWEFGBXQCYp0CDDzq8ULKO3rJdd8dER0N
PG71U1QNugDr0ZHQ2c+MM6+PolLEojIhQ6UbtRFUytKglM0RAB0cxs4h4w36BQzWbjzmwFIjcBnX
mr6YlJa2VwPdHjZfqi2q7fXbSROUtWB3agSJ4WSV8ULJxMQhsa28n7tLtQUY2oPwZnbOmCtrfmp+
0Bfs5EAD1cz2SNqjcPbsPRLGKPtMK6Ao2LoCr4FnROcdfM1wFy89pc2aua5FJMQqzSBYzXy/yXSx
WIG0FABiYD+5PY4ydUwo1RCtAFffF2DfXitOcuTOngqFj4aosWySm+gGDZ/ATeDIjz/jCzB7g3el
ccNDvo+4/VA0vnnaS4KRNpmVJnJbOszThSOKo8YokbRmDOWJH/QhfB6JfhQK4jIVO7IU3Cq/L4sT
LPtYe5d8wIDELOMsiFy9YMuZXMLF8rcUWO7q9EDEA3VXRdCZpKgbeBysjTxcBlrNsH3Fz2fzbwhV
Eb154VcFgJz0Dc8SDmLYgslY84/KB2fB/2/0IVZeaGkLQDptgXMeSv4XK6to0mvfvtd5IYAja6vK
ItJImcFj3OU4uKFzrkMMDrIlNmKvyykMHtDVAYeNodbaxqUsH9qUz5FhmSB3wpcDOLCBKwwCHCGO
8Fy3scewF/uEzZV6ICI0C1Ht0i6HO+77/AfsGjpbk3gzVUBNcNIMdiJzSZwQwnrF0L7Zwz+FJl4R
pUjsE3Iyn/uWh7ecvbS5RA7FqMT7LFv9JiWwBBqznrQ1MCYOlVDOYvo3Qck3vZ02pIrz18eN8TGu
KNR/HBYC4dTjeXuJzv14XgTFvYo1YF4HAgUbZ3OUEeRIjd5EAdiw1/d9Gju33QkGwG8BXHV/zeA9
9FZzJCT7G7Bx8mZD3Fo4dEBH3ZhZsKviEjng+0CKRAQ/5wiRkqsv/LuBvhP/4FGp0hOtDx1vlPVI
lEZwC6q3oCJLX1S8sEL4aGSK80XHopQS/3tHPezsg+dzR6FyPH3f9vySNhz1fMG2FF+Jp2Y22p1u
FsDRJANoBzYBl4tLfOe6lqdYeos4vTe1XY5BRxk5eRZXVAqdQxc3iVrs9AVMdYVxbc8L6QNh97sD
mQV9shB7vecSyqUZgjqNA/tWtkEI0o2RKkXNUcu8cvDsmH22yQHiPjgcd7X69ZRvTlP8ERJ78f0e
7EtLQ8Eiyq4wJfuVSE5Bh4JMubyQvkFd7VT7TtjrQ2+nUwDxcV15F1SWLrWyIGAyAchQ0cWl+Ns1
m6+U4BxoM7yx8yCgygiRW3NziJBWUvL3x6ZYp873GsHKND/ifkSFtDfmXIcaXwDwaHT4naQULB0o
ZAdh9mVYkBFLGNt5C5SChMnI8XZx1KGUwo7Vr8IkrrpvweIAOhlVt3FvfvtPIKM0hZOsY2apHE81
GPZsvvMVWQzl171lIynm2VTX4veo49/jU55sl6dXqM9ronjKOC/PNScYpaoaXVs51FrcwQgHFO8O
m8YQuOFER+8ouiXYMDSGZzBE3qK1KZmR7HDBf0tin9G+m+YIiYfl3WyP08+20ShH+3DNd4CWLh9R
89nlXxWhoGvZKt+4mn2JSnc/PW7sUs9B5vrOpMP04+wSx6s3pQiqqKgoTscry8PkePV5OJ7jygdB
CHrQh31QCim+WKT+Lyonnh1hxskB58MNs6RPuxIbXHVOWslIDkDbnewjAljCylYVXQBPUdW7IAsS
tp4t62kjKRWGrwXId5Ap6r0QMPROEMK5b6XxHyHp79YGVnicJCORaPsKwtHXRlAvbQGTeD2flloH
Q2YQVLdzT/zsKQnkaqSFjanszNcSVbI/d2Z37P7lfgTuIJ0cPTSf+EOBKQmyAVZ4W/WmTh1JkxbN
odSKI4r9X/UDwgvVO5bKxBI2tnmAkvNnY7y+ixKocHPQa6n5ws0v/snmf2vm1ocY8wnURDRLIP8T
WVno73KrRfWawTwtaiPGGId8X35ZZZr4OD1ZqJAj3XqmaBG36g2B8/0qsOLo7gw1Ni0nO3/2fmlI
kdzjto5V7deEyZrvUGNhmHP5FPLtzwKjICQMowcC/TW5sl9Ci7ZQj8o2VtZsGcbsOlkpgC3qBV0R
2vtvaPSWyk4dNJEiYOa/aofH9htYd3BldLIFOrjarAZLTAKeMfnt+CPBcoq+HpRRa8yXO5La0o+c
K9SJj2+Y8vLtdFwhhQKCcG1029UzqUD4IQ98jQZA7470fUeoITRIiN3VzDU+J0+3NIy5gTYkKTag
Hb1e9nz99wTgeX8LsUQWskc1SK8b0/oS9WuvLSQWPUajxQyo9XycB5c1HRTSbMgR2BKjt+YfPxvL
FGZPpzlGh670AfUuyjiBBAuc1ORqM6Zq4x2e2XWTrLgokm/dm4fCYYSScRxryyFTRGnZFShaDPH1
gphADp2S3tMnSdtfgRTw4XDJuMdkQGa6wLJGCy/6okhzEsTLzQcAXV2tAZIAd05oHUFMX86EoiNN
RJTIA/JdU9F0Dd/JrzgFp9Tg1JXZcAHYQEzdiaakbKgH/+/6+6Ob0VGJx//GLvSRv0HVThLxtmNO
DDC1NRFf2tme0/pyydUww52oypSVXH5qbacZDuGG3H+li+075/fczkkyaaCac6FPhX6FBM0xvn9C
PBQz0xjOFAUMLTIcsrWaGAqVh7DRpVpxFxFA0Glfsg8cC7SirtRL5wdoSKuy7h+Sr8Wvpnli3BlQ
GHK7WaXVcHArtFiIS9uuQ3ELVsJuZc+QEeCNcATn1ceEyOV++3qdHG6EsiwFtjK1t7bIDs32vv9z
YiDWxvmh+7L4/TCx5XnX69IZu9lejPuWnBjJdRiK1EKdfU5xgIcThbPQPHfF1wsE3TAYio7gvL4I
29M1BYbkrCuFfuQJCOfcsWYTXVAvlhRfXpXcxDtFxKhHFnN3zGE+HOdhHWBbSoOpdoe78dFXl5ZJ
U94WkStHR4zUwfh6NSQ77TrRmUAiaeuWZGRZDv8jJkhpdUF+klGaaMbbNC+MFJ9OM9BPMRWmPYP4
cKAbEd4fGlX9obQgG87bDRw0IjMIzaiYysRMjg0r3wMlxX4r5anYeXhq7ahHClivh5w5g7VTys5q
h5a8lg/xJjVEwL/W0rJ97mYZMYGYvEvrqoNHP7yOHobzDnd7LppbWTlO6vIw/3rhZSOTroSqgS8w
e0lk6JGWUqVK/0ZetYDvPzWt50huvz1w63KTZm1z1zKxtHt/2iCmrFodNy0s5AjL5C/1mHe2LMi/
/+k+zBCAyN0S7k1VqPvuP7ZQByDKWh8Mef0DrCN4HCgkNDLthPAA5GjDZ/+bKjXgd7LONCgw0Hh7
NnMSyJ3Ni/hYgiB1w1s3AtX4/BS3kWl7E77Mr1AzeuggxLbO5evHWgYeGp4mzsTKZfnJOX5zce5x
gtEi5Hjt1luDECPiHsBXMS4KRKwe5sUYyZfDw5GrR6kwILqWb96evTLY8a52cpqHUodEkwo2dItq
1+Japk+YL5gsGwYE9zz5EFF0Soaf+N1RTmC7fIEqnhFRlewx2rwRA2Hun9b+98gHVma5rW80gMnP
GGRtJMdtN3FkQNronFAgRNseHrjV2U2CGH/b/JLh8/Rvu15ov97O+6xah93hbJ992GfG3sFfDbzp
w6RhJGDZjtP0VOoOSrOeaKyLo9b24rIULLGLNCWjiBgVdkVjQu4WlVq7hv1n+ycixzC3+fu0BXQF
1k/aYX/5ciRweOX89Y03HYz+nc0qXXIxMJMM/htaa0RLyPzypC5kyLujXppi4ay3YKx3Esr523LW
4W27UD90ow9oyTufZ62G5L1hznZxBeLM3zWNtgPAe5+6goZwBDORKjV+6NfP5mcx8wrEK/yA/L1z
56UjFhp+dZogvp0MtQcmVqQwfjDoVE8KyOrpiFygLocgzVtPSsQtV2bOx19CiMBXFDbW/FbqC1kb
xAElSW1M5JZQFfiHtXOxMNu4HDN1JsccX62SCw7OTSNkXb6Byk/HNIVwamsQBTrjks9m5iXn+l5V
Eljo9kSpubS3D8ed6dt3/q4JOaE0WV9wO2fsZsgOzlEF50s4TqZtR5Elg+tWQOqJNFJR4xFcwatx
LDecNBGoInz0CQ1whZvUwAN8x1qURG7P7M0csX15RmBUCHS7zqalMmojKyWh/28Y7gsMQMfMq7e+
au+yZeKcH4WT+ecvU89zDgtCuRhK66LmPmvEFaZPj4e4tt/1ka4Tk02sJqPAsct8R6ybMdMRhoXu
G2SN524M70NXJMxhd+r11U2G1ezOzzOBbhojDjbEonTAR/wVvj3ptdRS27s5sXD4mGZj3yk1XoLF
1v2HzwyRD8FXSg/yJdk57il9KZTjt9E73Zc7hFCJyfJ1B6PDD1z+LH8wrXc0Knnf756Eu/mxouGX
KWFxrt7+0YZfpl++qAWsjHVXulCZ+4fXFPp1aFL3KG6cUnUH1sykYjzjdSYiS//jTMdPr6+pWuxn
vMIm/cevAYPycuonYTLzM9g6CrOD+WPvEk/c0BtDAJrhbryp9+YbsMxyJakCWSzqeJ2JJM4blZ8N
TV5pEntL3+bi2pDN8cgXAPQ/7yYrj85zq2O6fWfEME5/KgVjM/SjtXH7c9P9O6lXa1F0pKRVfC9m
kpCb4zRhi8YS7Fafk9ShHVXBe8VWytUooEtzeSOguenc89Wo7JnmB35FzKe4/THH27p5c05H4N7G
LZnExL0qzZWPyZXaMu8LupXEGgR9wrNtbQDkC6AlVqs5vdc8D9XHGp4+eWmc724X2Anp+c9tw5XP
d6MJxP/M8ec/ARbdq2LZDBZeDPF5J+4bbGar9S24f4pYZ178yMN+WgPHZ9JyyoOaFjhgGkwcrTdn
EBjcPc/iA0Ns7DFCYBUhBHsuX0X6rb3FFftY2pBAOP3VWse14ZWmIFXaCuaUO/8SWqZwQzPulb2H
5ocERTwMRRfBEFuIBxp/3V6IEaBEMDoTIylaPzQvTrwNsGFw5OSu9kbF4mQ0J8oX8spqaqFh8CR9
oYb9ShPY8MT9RvTLoQ9tQkZXXjV2YvjIoKFErRxb1XIoGwskUYc9i9Sd23KwYwP4ftcSiGaPe5is
aidjhw0xjY75W+jTDjBUwR2UY8EPyZWbbDbLOPn+87/bZzhS7cyzWNHZHeUmmv56VCelUIh94pvw
TMZsWKOMsjxWnV+oh1OSnj7fWUy2IrBEGCnXiWmQQ0BXyFgcfBKS1q0RXZLtDi+MPPQ6aB7N+LYA
z+GyWA8fatjQ+m3N7KE5P62PyR/t/KHt91SbBZKzpTMEztpJK5EXCjfFKTGHZeQL16utam3SBGx+
wK3Qij/hRdS/Xf7uW52bo9FYq4xM3ujEvcz0IfVuclA53Q85B6RCIC3Br8WOsrnDYTcLZ8IOhw2e
GmumjAjYlrebaXqmW5Z6/EcAeiwncoyy2O7RB6zJ409Vo6UpsvdBrlnt6UXXbGH3SidinbH1zbLy
WBOBOIwkvD/TgM9teJ/afPY6qhjdjFbUI6HGLn72nEki2UMND2zQV1BTLjBOIzRE/NAU/fFM7bb1
/pIap8lwI9GmPDZIJ07kR5aVxOcbbVfznZvfNF8XaPQ4wKUyaVA+rO+i82EUyXJo/FBDXorzpPdq
f6Vi1mHc00jM5ExwNZgpY44MhtgtNwaDscbGi6buCihfatBdqYLP2MZr7pgwaZHami7eqUYlJBZw
FN3Njp1+9qruGdCpAbTIPBxQ2udFfWBBQRqQrA3BNbdI+pqpmjE+59uPK79IF7NjaxiPWvHrq3U3
MF2FtsT1kFJAhIwEwF5ddEJEDPk9UrJm3qyeqDDDvOexJe9wfvbVtTBqz/stRcykxP+vfqqq4zSH
kaMlMOUCefBOsbbA1RM3IiGcrzAnpiDFgzu4o5Ma+QM7mD7wciPkjdQw5cp7dZJh1BrAbFxd9IbG
vM6PzscOXt9kFI5MwzXLaY1/8t9e2ClTsxT6l9kWn4L4ECSh7tOp/diKWFqvcWs4nyAR3MEmBPbw
g9qyXNwdXOmNNlNrFj1g36KFDkU1IDFx9p+8jUih6wJwqIL3m5j7JTx+KjnMZMAVRz2miZ7NqNxZ
z9zXjburCkzhinCkAMc4oL9uh+NQefSiVnRu6BhYPMrGW/qU5uJWZETc5NtTQPW41SqD1BN6PNri
8l39DKmmElYcR5utmylTlmHFGTrnXWU3Hk+kkLJXQzC2Wksehug6OrC0nW5j27j/1lY+M5mCwMrX
TDlNKGmWqiOd1Uc9OzeeSSqOYx6YtoZrlfiQ3kV7v1mPAFdKuAwD2ujGwc8pD9rFlc0OYw5GX9i5
5ygMq0tft78WHu46uazYmLyuYk+vWS96QZhvkIfH+09kpXo/vSIp7ORvu3CKe37bUK1W/EfazXuv
DdxrRfoBKbreeiN8RnTaZaYPO+IS0UeXITm/iGmAneTw2nuf02HUlNC9AWwTZR5WVCaBRXKsBGET
lqcRrD+5l+2cfKeLQsMmK71RMZb471uGUKpMr/zqKMlHVOD8Kv8YH9abziPiyO36GeUOSNQH6GS6
Ti1KIPEPb1nOuTjyDkCsL2Kx+hyGxqiXwQKtqV6jhb2z4x4U36zE6T9gtzqM/CroloeXCZvmKKVu
Jca9n8sbXPQMAfc+slDLPvoCBw0kiitCj0Yvw4HXkh2PnMBbRV25eGVVoIGLoMxXXGwcZMxR80td
lPJOYixUbUR0278Msv9DMgLwvY7FLH1ON7eaNVswTDXf+gg6fsXIlN4UjJ3F2uyPFtclwnQvjOxW
ohKVUNVxrIPjLfIDtMSIoBbJOOEJJTF3JbKxNwQ8GWkcwG8VJD1cQsJwLn/BrTN5sE64IS4Fvi/N
JtQYg0+gjIYOjSBdq5I1r6Re5SnAhdcHeSaljSVGBITFxWXi6ot5sahscq06C2UnhUaMDfUXJ+s7
bquvLaZkXMm/uB2LPLHv68KR+QlT/wNXWw4zWuzds+dmR4oVz1S9ZV0raN1wUWDDc7iVqNwqDkTk
`protect end_protected
