-- (C) 2001-2021 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 21.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
yRGT4lyJ0Beloh383Zg48QWA5Valk2+fj1pmz6tOGzuiL8sMlHPgB5GrFZl1wp0zCCQRlfmr8O/W
bfJWN5y8TIPAFLO9IoQTJIxePobya7INFnvXkxfFcRM2La8Xr5dnfaPVa6xDYaqIpXWUTfmwPF3T
MLUwTpctzKugg0TGwMoUlSdrzAisID527exn70nT1Ya33JeWFVmsI/X/wQrmgkY0RL+xx9/Xj2fZ
1GoiLY00FrRL0/sDx1VgscsGk6DH4/lAcKdpvpUpMvCc5TxA3YKYMo0iZVMpmAS8AOZT0bk635ln
MkkHIYaxz/qNrmzFjmc8FwKo8u4ysgrdfEAjxw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10336)
`protect data_block
gXvKs6QIPGqxmLhMn9nxQcF8z/3kW1uU8f56e4q/NGV7Adj/BDrZ42h/bfTiLcgFv+GEPL4MSsQs
n/tWLkldLJrugoj2ITz40D4ltVoapVFCBkKX/6vjCRGACOAIQNwvfhM9j7/ifBMLDTO08V0uxR+E
BJoKkXVXXZFvC+0vhfCgLmUAHaBB6bUFef4HBlUGVFiEcRjNAJKrEZoPcz1DiBs9OkEEeA0sVs1p
ByEGKZp1i6VxkAUSsaRRyU34YYPjlDYLfRPMlmO8Sk/XizR2tj3JUZ0GZ/z/NU/thSJhpyvGO2fj
U53eCTJxBAgq7sboeYDcSuAwfDPQWkm2sr4HpN3i+H3p/10C22iRVRSQRxMWpVnNTKIY+JqSmcGK
FjV5BPdFX59CFvd/xUegmI5G8knmQeSR5CdJBJxM4PAq62zcxfCS4IThICZTOkJtpYUYIR4UdR7o
9+wBNw/5MJXLybCuDko7j4/nXnM5kYGJwE62n17TqFN1NS9QZ34IQiKuMnrQfPUGE8qLTdzYiCm6
ZAy6+ztkIDtENlxfu6ZXRqNDSQOvcDnCs5Lf2uvsfdo39kXTgpQkpnbD7j5PzqZfTezPdLFOTy1c
23Mijdkf78o5EpMSyx35q3zwhyaYA7D+uGkxSDQsuQewsLD4cdjsTJdiQKpcQ8U3uTUVdbDFTvTC
SNW5NON2XEnQlTI59wjlyS6phivD53/oda91KZFMMcqmm0uTzIrddu9Ls+2wjUrm4/wu24vTuvSZ
L/eNxhY9wLKy3JGllx0rW0pAC//t88tWK71sxNMmQ5SxlMhnUR7rhs6KdKYKk+pmk/S+8ujqDWA6
ThdlaPLcwyrU2mLX7xYT/it8CI1u0FYNdVXjH6F/pQsg1MuKFQ0soa8XZ1dlyTjdWGOOc4bsC2Da
QuYAChPD6l0V+pOdlFdlHkqL2MeO3NemIIRlD9CrWTHpGzD/y3a7llR1q+xbkTe5OU7SWzEp5o7i
dFi25Cdd/X+A5glxW0MgWP5M8ovF5f0mLOyHMRrr2R5lUkuFHH+tjY01WMFz4xd0sJS+qRb1cIDG
7fJmlCU69QYX7JY4owhNmKqXF8o2pYc3B78OnL7BtSy3YyaFyfPb/u4pygkF6xsIUu0TiJtjMJja
JttsWudhpiGm8weZ6JdiV7AIKmq4Qoy5bet/OHi4Jf0N6YLNJDHnjdrn6VTnGnukIZUlUwJiAhQA
kyA2JzNhdXU5nzymggIMiOfB1KsJROJH2rlgAyZNGGOPVUMNdfZj1tc6hIyCMGNT/KWbnIYQgdgF
Cg9c9Q0A7BX60iPekvSPhBBByphKEL57xywACaZv7m2Fb7nKrKt2+dUAhxyZMVDPp7dAe17zev9Q
KEdv2Gz5SUa1nF4RMy/Vv+zildy6HOXpmCR2+IOoqE9jcNSEbhEN9Ti67MZVVnySZI3bxnOkP4WK
kOC9djhhApDXij2gPVi3yq8oA1QrbNaYJf7cpRdHwCUvu9D4o7wZW2JXa/pO8SEt3jNSq5kDOj+L
pULHf2Epcs3njXqA5v4IUpfVEiG2jNOEKk4S/YfTqM7WpqlPBsAy2QzrGM5do5Hr8qmkCQqkg+fm
dfwHFKnZs0s0UJ+mr68tyaZwg1Mc/VamW1kZBBkeFC8aV2ImZuUxsc2G9Q25mgeWqtcu1bHQBbSk
ItP8qJWHokAD0bKRFgZmguYAL4cfz/fc2QJdpqaYkjPoZvp/4qdeTz1CgQFcnJAx4mQPFumquQ8S
p/zTD2QCIGXD2up3EuuZngNef6Odj3T0+kZKmwAakvwTu0ZN2xNsxOftR+h9mAwpdK3Sd5hzmN86
Fs7wcUFhklPoihCbcYrsveq7IgV1tdNtzLydwWe++Pr/luy9wkpFmy/dhnYd3uldVY7UiN2JCH+O
EPLNILggUQ2gSgkAO3wWEfA0bL+sVripQn6FXUzsVe3XN0GzYqEie0Qzm2Xu+pDfd/D1GK5RguUW
/WozK6DoFuwVfo4aFYPvhl25E3SEOVovKnHNtww110O7CUx4fOCF6kRXFKMkApFacTyavgGT1QIs
+hpsC4mfmHq6Yeeh6tm5+yHaiP5O/eZVl7EHw6GTryzEVi5hU+q5xsd1iuLmGQtDvjCqUlWP27LW
4ELx/+u8FxAwcQeJEqJJgV+xQv/eX0hsJc39VuqDc3Wx+d2COlz4VDhUr191pCzKtwcgLlX1aFQJ
6skAa9ssysNjB9qmbOgkuPiY55pTfTh0mNU8FP+/FqT1cuxrtBxYXsEzbN2Kiqk/jBnd0C3gzcb0
cG8jy2gKO0+PhOZWUTz5DrI8fpfxYWi7s6rWPOXURxucjc495o9zPk8Yo80Fx3+k8QwkI1P3j3SU
DKfXraocC4A5T5m4Grlh20qgkYEhV0+TowCb5XIdXMkZjx6FEBIabmSVA7Cu2e4XWZIBI+dNgl66
weWakdI9MgQPcpjKDKEI5T/w7HupmiPbjLK0st/CPDMbhpWdX8q9R2oI/gOCdMEuOf/PUA0eikuK
g0Vv0LwTZ1511bD5PYT9RQ5KRYzUeJuPBI4M9WA69FDg1Kw/NJHD5+BGP0NvCqJeCcV6dNoh/8D9
TS5IGbKio2QKOEaSvQmyYusa10XI9FRIe/wM65XJUtm0oUosk/mBL+yIhTeoJPET60Ee9P61u46x
KGhc3tfjoO/KTicAeejTK4RvG+RxLHxi/aKuJu3Nf2a6BdmqjZRSfYzldHW3LaNPX9J9SNbmyn0Y
BHO68oceRyjacdK8pqjJMcQKMZz0teTZDY9jG7gIG7HTybOixaPZe8zH6uMiGnE9bueSF2oqGMOG
1uRIaytSJPxKB/iE/f0SjQZzrG6dvwjwvPW11P/t5VnGeX0i4AeUQ+aGPUbi8JEFnpeyV+koeYjc
qasdiiByPGcpbueLqgY+ob37qlsAB2qsM/w3t0BY01INf+U2tvEoVKqfskTu0Vxs5mmx1jFvLFTz
YEVzv5LRw3hWzOSro4RpjSphzFt5Um6AMNEMw7/31U2YJaWBGLVWLVNvjG73lh8X/7wV2i+VzKZ0
7dWz0MjyOkK65psSWaKMoIrJR7kY3piqLqXMnndytG1xo4w2rdl4Gx3BJHDeFlF4fpQ2DJ3jdAv+
u7TNd4oqCLJDSh6d039B+5oie3Kz/MYdeT2J94uzZwbL11sSbH/ttAMb+4D1Nf2RBpNCUwqKc9Q1
fqmoRZGksSNdUkUQA8zWZCIT0zj3Ynk1evPisQnrARcVJfS/hEmwgRSaEyRhhSND9DdItm4fVaa0
yX4dqWLe1lk0ceSlImj5IOetGZhFHx+Op/44PvCESkMBxVWgL43/9RGiKsNlBeId0oR7vM04RvJX
joGXc9VURVEXOBx8wotpEyGnNgK2GRRog2leOV6FsclywVGzxPe6c1GzNO/W61akA8couxyixlH2
LIDozl7LPKRRT2QAyRFfe7ss0UAV+fPNynNe73TgRCtwbP0lfETdimwPwMvGiqg1r93o8vr1qGkA
XcTK6qwtEVmvyms7IPs7tIttq8h7hpiaYTmbZcw7BOw3/hT3i/7YV9bwXx7fbaWBzh8YxKV8pLBW
4IUoL3N7R0C3zAH4RV5y167mF0dHSinH+bv+1ckzVkzSVY6IFkbeoYkOi98ROwbHIy3/xxU8XS7e
0Z65WZ2SSIFyxUklfiRVvecoVzKS6nHzcGdXGH9P5U+qXF8GGXi9pXJ87h2MpR8mJ2cM9vOguTmd
yGLLUDvtEDoJx99u6tqP2YxaCsVX4LKiOfdqYdJgGv4px8/+vxVRYoW0GfqA89yC0uQ6GoFwdl3a
nQ//1NmUJpJmnmZ+smxgmx9PPo1p1gSwQQ8IVzF2zUKUJSagNJvQKvJRjmMpdg3grxULvHgLYV4c
K1gscxLEzTLhELfE56mfsjWb/NA196tdMdXcmv/IkvV2MOvCqiOyX/TAi9jJiXgUHr+xW76Os/01
oscvkQf9lGeHvidl0o5wHJM+3wqgk6WwHAPTrIKFmqF6/gqmJifc8xDl2hMJkwiBrCKpZuIgL0in
f4aCvL6SdlOQx2K/5jq7LsaqZB02YopBhakk3ZKnhYENbyqEX3JpKObt6ULxj17nI15EGtcfylKA
VO/kB9AK1hgKpo9+ND4izONrZtM1IHDDp/Yddkl3GpUh3T+c/0NW7qVysGyxTdy5xXOb/p1cjAlD
pjV0/a29C8YGbFBqbefO0UO/nIfP9ctQZRRc2h8rOxA4FDBFoEuEJ98Fru0FeSu+OCcYo6VRqkvu
bGng2urdaZ1q2I115FHfbs40rT9Iyd50PTELwjSACB/Xemm5kLjYVhq4UOzDilf/fc0BggKBgT5s
wMfMuY3Pn+o/xs9Y7fB6vw2YP2fQthE4rjDsUE/WfzFl+EFixGSKW+31z9+kEVhoTBwg9snH6dbF
npBXCy3tvCFJpZHoXR2tmoIQtFBpwaB3vk9hSsUJADUJPULsRS3wj0e+LRpPT3FUayzqxyBUvAY2
tKBmm1oBazTHPNQqH8VANVRQvsQzLzIHejDhyv7oKlvj4bS4z+tbW481Vm1BpETxFBh91E1Sub/W
WMCos9smFx7D4bMBideY+ILQbu/K7ByyB1W0rlIONUJQ/UkZVluNR6XBLTp8W2SZ2ViLfBVAarNX
oOQFWjV0wNIq4qfF0CoqECfazMuqc/irNLsJS7q7rf2Wni2TRw8QveoH+v+Jpm2H0ff5jpKBcHax
QcxLVZnRLqkAvYNC/EPIUzaaGInES27CE6JbkEolnxWSzRJotANy24sedj+lj2kYn5PKAorZBYe/
TyhfkKMG2xn7GjK8gKpB4puW+ceMWPILtLKTsNWGxKFR2lRHkGxKcDsnO40DRxszNlxuuMio14G5
J8LCLoe/otGtxHvwyIcsU78UXSYWy7WFirGUY6Xp5CKJApIzm140wrgBJCy067akSTGFhefdLbBK
2k1FCr0O2PTCJ48XUebU5LisUzBsSKADX0u0pJWs+jP1/4DSPtZW4wBJCgmJKCigTrxlpRa5RqEW
mQa2wjv8wVzpb9ayksDb7VB4JjYdvYtt107psuoAWOns1qQh1XlNOr5hhhkNi2KOW/VUaOs813Gb
+fGMY8fHjWgjgYE8EAqCr8Fm4HpLVOXQP4BIRQASHCExAYGIpCQf4H+cF2Jnrdv6Nz9P6BrPgjZz
KfHXak1a7+VbfkxXJmH2NrfIwtm5Ll51wCIWwCOe57Jd0N3P2SuAyYCAW2kkphyqOkVmZAJrxY4V
ujjsom8WB/+GnsvattkUZyfNnd18MlFPFZrQbuoSc605Nzl0WpFvyBsw5GTlHpze6d3SpBec6J8c
7v8/sEZ/S/GL/Y7UKhsvkP4LQsHiMM5lCDEfisAjt0KD+aRaCG6xk5RSV/Ch5sRprHx/D7O3WeQT
6haT1O+gJ/eaOj5bN9sVKdX/sIzbzMxd/BKlhkSyTATGGx1TjOWWO62q/N6JzcYS8RcCGrwpyMS5
1rWPLTFv8zJST9LdCPkcS4vi1e3/N4GNfWPj6D7QM7h2VcOZaIrfR/GGqS8iC+wz49b3qeCbSB/n
u9tEDq5rkWcHfRexstosxIdSNNkx6PrpaKULK6a3zndYrG4QEHr8zMJsNNDXdof1S2v/njHonR7s
af6PKhR6iTthyndXEF+9WjpM4M+RGxzaxKIW5OnL95N/6kbTDrHPDM97E2qrv06q6AyK3SdgBWt2
Mn7LC59SMUkwl6LSpYlSVgfXzhusVkcZziHwCkFOuM+yzzJjgwv87GBQV/W+SB8N7BG1+7SAeAC4
lblxgHGb77qi/GtT7w6gMxpu3B+Ee9EUCbVjHbz3CLwVWZf+i/hAqcKk/mJ8fbJF3382VyYndhKb
S950oF5MRF+iISgk+awhviGj30IKZKWta+NZ+HGmJspJCad85uBHpfSQ3oaxrrnaXyJ9VmiS26+U
90Q3Jj2E1fY2S5/GU8OhqLWqOY7aBvooLw5xXWlnonTsUj5IjjpD0VRqbKPha/gVRdlG0I/85+WC
Wc/E+Tq8lWH2jAgIcKuPXvIEzB6ue1P/ibOWf96I/cgfXUzpsEidJa6ESikirG5ImkxDfvWh5Vx3
E6uocW+xzxPmpBkXqEObC7yA5X/n+RdoqityKI6/2AKKhxlw33ZOYy8iL0Q++2tUVpr/aE5ln+ad
QWr51ZVZuEbPBvvHmGjAOQFbcrHe0n4RIFJeohx5UO9RUn2B78nrGQfjTtqQJqoK400f3MBzGrUk
pA4HpWFMhsWh8LBYlDmv2wUk0SiQAxxnFEvYiZ9VqWbSYXoltWMFpd9Cny5B2w6GpbuZ2XT1zLu/
alFhJ2DVaouhsawEJ3JI1ekAdAWxz79gNfVClN5sTqpgkM8bZ2VnzTO1TAHYJdqC7t6OlSehzJSP
HZ3WYRvyOwi0MSk7zO8Z9f16VukjrQvw/Dtd2/iZQsja2jwrOz0lpIaNiLjAstWp2k03duhGPg0M
yaZ4FLwHR1x5msRrxJhf4CBhiNe6uZFabtyr5AZHLwNy6NA8t4wFVzd4VD+3V8UKtfZqMzmVE8Dg
oqeTXCp3yq0/SHpqoT3Hxn2SVGIRK7YbzEkq6t/yI0UpY881Aygq/l0LVSHI3BPRIH7uHVAA/Ier
njzcFktflhh209nF7ggquittb3AENkOzW/6VptaX10e2TAosfrYH0BECaNJ9v/kNMk317ZTSIRr3
2D/0draDhNRJmiQNXkdcZ5QNnvXuZ6tdaD/7w7eneW9Fau9LnmxQMyekkUFdHPscdUueSvYKNDcB
mt/DoJfJc0frQYZw2TLiFMRwWvDDR2lfDDaFvVbLdX09xXIVuCi4+B+wtr6FOdD3ucgu4C2LdMWa
3tIcRAk5ZCA1CgI7Upxm3mt3vjfzukBZrW/Vy436/vH7sp8GbyBoTBmagNCiJLwWziluVd+2xrI9
9AncAGa54I1E3YBLdIlRekxi5vhlbUvjGR210blWVeLaaf3BceAK0vrfWpLFpTQ5GeiQQGHi7Tu4
znhIf02n9wvq3+Omu3ZtFXF9lQDq/9ZpdggB4vRcnke5M7SB7vBkdPD6OIy6NdtooRc46wrExU4L
kRn204eT0mqNBHRwgIFnY9y8bMEZY/bYk5KpEfjwJdbOh3FVbIqTP/gu+tZtXNStetmFWvy92H97
vtLizW4JUIiQ5ubH7XAzDAud93t4xlv2ljshLR0oGiPGv5ZKpjV83GL88qW1P3tC0goQihn2h4TU
O4rXdHjNvsL0dNDGf/FiYhrS5RCJAUPppICHuhewDx/ghS2VWMev52Ne9ySkkU8G7JGeSQ586kV6
YfkQPnBwH/0bw84I+nnlumq0sqLzRy7MZN1xqKnsx2iyczODLZm8YKLSWqtZK9/ypX/fyfj2ok4C
lCu3fYkUqRfKCW61BBE8SJIKZT6uGZYCOjUC78kqM2tpH7By6IyvBrcllDvaipDx52XPvXrPrYUw
1Bdcaaw1zyqcVa/x9UjsS6xfmn9zDFgVrgKvcaHH2GoH9emVYeXXN9HYO0bfnQahiQU/YQVSgi1y
3dlDQ3PAuA6dMQemxuvQb7kexUyRiXUbRHPqGDASXxBPRmbfTGUYUizYtHXsBroaqBHyNCmk3afu
RD/EvoQsSxtd8Z/hA945U1oXePPdoSfZZgpbOWDfzce9OFKEo5fAJVpmVrP/faA2M6lHItm5z4es
VINnM3654pUCUBJHLm3T5sl97cgj6rbdGkEZpA26172sB6zdcondLhJb6+oqeK6VsfSz3oXNU4KT
+MKP/IfFPPPIYqxWXmRzMUA+mKVbAUVmZB6iiA4sSUw325YQd3ej00duwqoabWSOEpoN4FnNerXa
xY9GeW37O1x639MhoQeNLuVpk0daNG2OWVSF0MC6RSrcc9hc4YpNqABlnMwh09jWN2mKHg/8bQS3
TjpxwI4YrjMmjegVBWEWZ8RMBiETYu9lhdgM6wuXHiPo7N+1efxzI5mtSlmgot5/AO7rVT6dLEG5
0MyfkUdywGKTT4G5tOLjPHSezAuby0HrWMT6MnFNFnKnwp87NmXEEXLd2o6Nhw9LWE3Zo5o2TWoe
zQbYJzy16i4mCZKI3n7QlFlISUVcc/V5Qs0b41rh7Xe4H0Jn+gh1uiq1ka4zDblOyRQPtEM61+aD
WKKHBch6lZPBNp0g0Wl/4SR5OlS0auiq5EicNcPnPctaMRN/Gos2RTHaxpFjdDBRQs4GaHwjK3mc
M7Jza3LYUHbRowZd79eBF8oV1mWFnEn/uoEZ+u/VB5vSEfSbDEt2EL8+iVv4QHjWl/vWbVMYoi2k
fClgYAcmng39n7If7rEib7VWcRPddqs5CQjzJH10GdrZVwEgL9YqcC1s28e1JG3uug93lPrDwwSn
0duTn3f+m/7tkdKt2e/02ww9Ch2nKUWIJVzXvGfZa7quxSKzhf8usWAzClY2JpS+1WzrpUPbyBzF
gf0i3EhOgEbkLlnEKiokVK88X1jWq4WtmJ6VJ6D+JGl5748O2/6ZK0+khlGrVx4YIiBifnDaGa4c
8kOH89sovFqAHGMRE9JQ3Vt8ldYemLBM1gNLOSJbSotclgviNJ7BqIzZVT90kDzut42VUvScr0zF
tJ4SI20nqRdlnS7ULIgcp0YvMJRs5AkLg2/oV9ryC2W3QkkUBC3MY6XcMk0qTP+Uccbp9K48yAqh
hjSG92UGJ+cZfWnQgNI2VlHZo6UJJcC5Qx7yLx34zPIIegACijXMb7/cc7KF74C099YWxtUEY/Hd
8BlTDOYfHHZL/RIk5Dwvg+XunwZoSHUZ+8qyNnQOmXM5B/hCUvmfajO6Y6NfHyVUJfxH+Rkgno3l
zTAOEyyRd/6mbgxagmHjbr1XuYEOGTTExSB9H5L8ldwkCJOcbg7L5hheMVUAuXv7p2asVoIAY4Pq
iibZkoxAKsnob8hqHQRNbXeIwBE6G57qvJPDTQK33iI8Jqv/8ZqNWMwNIws/vh48p+OPkkhPQatb
CqxM7ko3awIIPEkp7O5N0JOktzfl+0cQX4Obf5v81a9E2bDvt+OGThYk7k2dIkLH9NaLRSOqN1YG
tXNaTmCFeWLAJfzxZP+etSYD62mhTTUpVG8hthbj/SFxk+xSEJoEhKoms7JJo9S0E9p5e0McNkMe
u5KBp7Ba0abwoihaGthIptBqL2HFnroeHYDXsbnM3r/aQ24lUE7FS/CLRzEw6DBfLmlZNvEJIAeQ
EWLRqPk6W9E3YMaADLV2DJHeY/KOQep1PhLs4mkyILoHy2gPwvnBawX9gSXtefk/TN3f0sEiyazS
Uz/EHBouj3fV2rYDnnb1srJctUqUn06CsIN3s7LwKymU6OrDOwqmRMlw4dmkTlh9m1IK2BquHYBU
d7fqdHoEEW4JB9D6zbnIylm7StV6yDc/Wj2Xy3XNA1s0lnSSZ7veyx1uIV/F7FjghLGdmfeZw/Ki
vGwHnTIqnLfZUlG/oU1qW93Aw+nSggG48+P9R/D/Q4TiaM4HSvEfJfBVacwi/suO4Ek+UFZ3hfac
wktwwkFGskAcKvnjlOhvTQXshWVw2MWAcfw9OFK8APJIKRnc6awDMsEx+yAOrZNPQxLbTboKfwWQ
BEvlkii3EY6+SwCIhpWfjlHj7N4rH7v4XHlj6DEx2cngNtl7ZYO4HjGoquftDdqVTy7zKRzBjUqn
dG277hKANOfJ6Nxda8gZv+fbs2AtnzPb72KugaXog9rAFU1WeLIAEdPvDE05MA0NwRU56LRl9f5C
lPtT6OLQ/zNX7FczDrrDDfLOapm/OJeaeID5NcFLXBRaD1fad22d/3XWbmSmNJXtuHWxK/eXlLob
W472J94Cl7w8Nc5w/9HhiDRHq9yFIUfyH7DjSUDpurb3WO8AENrolGrE4R1odvMhERkf+GYMAI5r
rS6rCP6Lze/qFwajZXwXrssZfxuiA2MA+wG05BX40BvXz5FMzwZ3hyV2slzboKo1DlmE9TvFxgoX
9bzCHYsWU3KPzq3pJTo+w5uQjIaCYLnZETYorMzjhAPo6a2t7+LSZukmRS4G758pQUxk7VCHtPYW
XERICrOe86Tl8+SbioaQ1ms0s+1qUEO6BW3b5G1qunWZPHmEIfDdkIfySVpuat3VIN2PFM5AkOBQ
Y6iG0OknKjSAZsWmgiOsebFVdsom+9F13r/gViSgWFuCqHoMUzDQbZO54ZXdAvbnq7C1S6rUpzzo
U4gl9jus4vHiXZkbIY5HmcDVCkuSsLFc9ER1esDUCZhcg6KMp3piT26Ck56bIzEjXYnLAih4P1aq
6XqzyuyTYXzlFiLlZLEQLQ9AiZUQcApy2INsLLGhU9fbZcGDy+UjbbH8AJ4W3n/v0oH5UBKbhz14
2NC6Czva1OD/W5cgp5MP7B3i3c3J82uoC4al1jSYvnyTmC9mec12IjVAcdyrZ3HcYxGlXweW6Arl
28nX0ZNxGqobmovgJJ9dybyiHPhG9LvjirsrAR9pQBc4tjE218Ousq/H7R2y2zRiB6NJr2faiDAB
8N9d5QNF+R6t+JQifj5cTUji0XQTP9IzGOsd3fi+g6jc8hOym00ddxtm2/VQ3VoWJ5DT5luonPWh
CxkmYwQIElRC+YmhhRlFD20DnqAGGAXSrGgu9wQdjmWjLTV3YuEwJ6FLAnM2HOu+G5N8j8iJO0Tg
FrKkutGaLz3JKDuFsXn840RkeS943TNACmLMS/89wzc+9anJF56rfhWKAX/ph24JMCV9pbQf9Jvm
C+oEuGWWLQhJ5JDJM/KLovteeHhkufveIoyJ5NjvavqMKB1UVL7d6vae2LrLn1w7toniFCBpo+fA
PO97kiN/L/mi0ba0To0tgjGgv90GyLiVxICBUXipU4I70/4pN+Rroj2hYeG8KUToVkuQJ7qXYD+Q
6ddmL+ILxg6bfFKJP9LXhv7UgCsAV5HWLKBP6Uv6MSbQvjXaMak0dVmctUM6VLkhJkYWiVGBlc5j
NjGfbxPnXuzBeErOQNAf5ZGQBK9TxrdwCzwqnbPx6G5gJVWx3nwEfmrTzolPNNddsVn7ddSRinD3
SI9d4Gb/iZDt8za0H3pyUtJPneguDNmYOFYryATDYN0MLgzrRlUjnimduoh0Jo0R06AVb6lPJotL
a2IAb3cAgYxzVs1BBzw9Wg3x4vs0GARx04CyxSCVac+IbqR/BQkPD2hbHgODyNBOFewnoUTZPVtw
Qs0JsFzO5ZtyPusqP32AQsg9HXQbAd0Rf0gZ8Swk1aA5Jda08X2mPHk4hy5F5y2zzbVf1qe6Tpu+
DbIps0WZZ8ycvFYSKqBVhilbs90LPjU9olid5Wg25/OxbWzDJoMBjtV2CFh6h5I3qQJOo6nChrF9
lGD4AZFzDAMCRb58p1SQ6eJi4fhTz4Mb6OMO2IBDv0/1QLEFBBiqk4pNlUSdUrnNZz9l6hyWwMkB
1Wxyw55Hdr53ssJHMJpEALWeAPtZNFdArOhFuXBZ2YTbot6T5Za2caCmoiAWQjnEMPbkVdUUHHtk
YQzyeGW1qyvxPKd4lIK8cgEeDDhxUukV0sp4bLfpnDYZai4HltwwEVkbpWAV6Y2dknzTYPrtw3/D
h0LD7A9uXMtRD8X+ZI8X5b7fFDtBl2EzxZD7u6NIY952DB/gzqi1uICGTi9QLuWN8zlkhprhDxzI
2yh7ZF6cBXN93rmba6u7PZb5Rq5KQvPKQy3hZIuakweBhaE4GXG7MQMDk53iTDH/WSTQyHf5ND5j
BihbKPTj0OgaU2ofGuYVWQ4Wrcivr6keQvwIYelDB9ZGPyh6ZPLIBmSRG3D4ftagEbhv/RAqXfl9
fiaLt6xjLQOHDqjgWqoP25ml1q2qvDmiZgTaci1QzYWxYNVTi/yKsoVcxP9DUwYyIE4VGjyxaDM2
TrZTzP54dc1x5qohZ4KLGgk0PHWoo2to/RyUiTo6x/eCQsX6AvIVnEqiCeTyh0oApO4PkzS3ZhYS
zRH44dE+ny6fQKVLku6Yut2Jnr6dCGBn4XlVZcf3veqaK2PL9NhXcx+iFrYjMtldV6ZAEK3tB66r
xECV6Pt1qrrDiivCA2ZwaMnSLJXxTitEAkbLF1pESCDiMP8vGyVcIEIT+azPuHGexgp9g5QC5B/z
G1axZLqzh+BGgbneJytOVqqgfFXe7mThfNNxj5qYR52uZiotL3tFgCSS8hQMXM61di0vD6SXeJko
eAuVN7GvWvd9ShIp/4tPbQE++AMG9Yn3VBu2o4J++nwM5zynzwp/Hvubu+D15RmpvLF1/cC70HEt
coBNyBYRs/+iwANvU49x76FwcNRLkU1Ro9Hc4Wi8iIm4tpekd8lRDumqB/Thd5EiOj524zcLZWZ1
/sLgRrWwQ9o3ZnEA/0ghfynCq7fD0FdIV2fn77Pn9SRxekXcVgB9JKT867w6BnSVIkpHBb2gvAaq
U7CT+1qV0tUWI61LOmNFc5O5aqQWy03wkQmI4oke5+40hJv3t2HgL7+Jd6XA/Xg9nzJUDei0pIlf
YvN3plCCZ8IIk98vEkwC8gAV511aTPLPI8BhdZUU8oQTEKFBjYfRCehk2up+b+6EfV12PxD5meo8
H78SzWkRLViC1VqA2R3VvvowW8O9cAdllzJ1lKx+CvBnrtdzG8TehOLRS4vkvD7zAFaZrp/f+B4r
VCMziE6f7aot2ukBgKYxc56pPPxQajrc7bPm+f8pvoelYfobTpIH6o+I/gwd1nEKotamakd85NrP
NdLNyGp5YESPgTfAbvm9W1KvzD8XdBXrcruOm1YHQg+ktEWesVPDHaKxAkFvY+PPRuWAPUBOIcTF
6m3QoHwJH1U+8R5OpGq/cfpVG7gFr92flOGfj+CuYEHxz9duLd1yBOo0xCw/lWgkI/+czSpDgRzz
Mz202CAjqmhHDGB65fyuNIwB4/4hYdkf25A7hWRCSRGS1lvu3KVyKR54AooaePwIRWKxLfp0b6g0
wJgfwzjCLJU5g7zfyxt0zQ2rR8O25xvkzZIrREL7gTKBNx5fhnSMVrXzitheK/l5Ps1YFCv/s/Al
IhcRJwNKvIoRSkNftidtAhjEQYlcfaTQ/EiFDB9QHBrtNE0jTcgfrWn0ZntcyHDq1cBPM2hYeQN8
lho03HvV/DUM58VPt3XnTh2dp4CXuaE3/5dz+LLMHhSq0I9k8FF2VSjUPDinPflPrSGziT4s+sHj
FaFSh7bS8htkUJ6vNoeOFCzkNkQWGvnrGqaZYXmtGPl1CCxDUb17ASXfyyboHEQjrPxfDy8czM+D
fu9Vufjcy3vT2P5rBtceQuWIqHlLKjjnwPYHszYrtoques9M0JHIlBHX/UUiHbsco3AECncwa1Xp
p9KRCBri3IncTFRz0KAZ0VT9oQPwXyPQFZsSacsKv7VIr50+xqIR5gOqdXNAT+eMoNTxKXyP78Eb
Ew3m50z0qPdTVlRB4htg99KOP0LStBu8DT7fW9ZI7fLoJH6IFuQnWQBOtGj6nyb3E66xNZDCYdvE
zyQGCfcQ0Yz2KUJwGZBEjayTE87esMcq5/zWfWtuNoCqSpWbelchjMNCC6aKXxF6gdsrQQEMTSAF
hyDzoAi/icwGBEWzQMvaoookVBaNfqDzqiGYAXwdvMhqQJR4vkS+9hA8pIhAm2HdhRHoD8Z6/w0b
Elk97YLpUTJpIS8SnU+CCQ/bTZmxmYVs1RYdvb26lkXliqbG7xBZWTzQyqIk67GOVTgNm6WasMu/
c+mLLJ1ERYYHjy7hr4EDz1+192Nnhw9nmGXQfBKswreo2PQ9i0byZZ1z7DVYgw2jCoL+7TSa0CWE
kfOi1h9I7WoJStczEErJELufpw==
`protect end_protected
